* NGSPICE file created from wrapped_tms1x00.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

.subckt wrapped_tms1x00 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] ram_addr[0] ram_addr[1] ram_addr[2] ram_addr[3] ram_addr[4]
+ ram_addr[5] ram_addr[6] ram_val_in[0] ram_val_in[1] ram_val_in[2] ram_val_in[3]
+ ram_val_out[0] ram_val_out[1] ram_val_out[2] ram_val_out[3] ram_we rom_addr[0] rom_addr[1]
+ rom_addr[2] rom_addr[3] rom_addr[4] rom_addr[5] rom_addr[6] rom_addr[7] rom_addr[8]
+ rom_csb rom_value[0] rom_value[10] rom_value[11] rom_value[12] rom_value[13] rom_value[14]
+ rom_value[15] rom_value[16] rom_value[17] rom_value[18] rom_value[19] rom_value[1]
+ rom_value[20] rom_value[21] rom_value[22] rom_value[23] rom_value[24] rom_value[25]
+ rom_value[26] rom_value[27] rom_value[28] rom_value[29] rom_value[2] rom_value[30]
+ rom_value[31] rom_value[3] rom_value[4] rom_value[5] rom_value[6] rom_value[7] rom_value[8]
+ rom_value[9] vccd1 vssd1 wb_clk_i wb_rom_adrb[0] wb_rom_adrb[1] wb_rom_adrb[2] wb_rom_adrb[3]
+ wb_rom_adrb[4] wb_rom_adrb[5] wb_rom_adrb[6] wb_rom_adrb[7] wb_rom_adrb[8] wb_rom_csb
+ wb_rom_val[0] wb_rom_val[10] wb_rom_val[11] wb_rom_val[12] wb_rom_val[13] wb_rom_val[14]
+ wb_rom_val[15] wb_rom_val[16] wb_rom_val[17] wb_rom_val[18] wb_rom_val[19] wb_rom_val[1]
+ wb_rom_val[20] wb_rom_val[21] wb_rom_val[22] wb_rom_val[23] wb_rom_val[24] wb_rom_val[25]
+ wb_rom_val[26] wb_rom_val[27] wb_rom_val[28] wb_rom_val[29] wb_rom_val[2] wb_rom_val[30]
+ wb_rom_val[31] wb_rom_val[3] wb_rom_val[4] wb_rom_val[5] wb_rom_val[6] wb_rom_val[7]
+ wb_rom_val[8] wb_rom_val[9] wb_rom_web wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i wbs_we_i
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05903_ _11560_/Q _06228_/A2 _09380_/A _11550_/Q _05902_/X vssd1 vssd1 vccd1 vccd1
+ _05903_/X sky130_fd_sc_hd__o221a_1
X_06883_ _10253_/Q _06883_/B _06883_/C vssd1 vssd1 vccd1 vccd1 _10253_/D sky130_fd_sc_hd__and3_1
X_09671_ _11633_/Q _09669_/Y _09670_/X vssd1 vssd1 vccd1 vccd1 _11633_/D sky130_fd_sc_hd__a21boi_1
XFILLER_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05834_ _11687_/Q _09998_/A _06924_/A _11734_/Q _06344_/C1 vssd1 vssd1 vccd1 vccd1
+ _05834_/X sky130_fd_sc_hd__o221a_1
X_08622_ _08793_/A _08622_/B vssd1 vssd1 vccd1 vccd1 _11165_/D sky130_fd_sc_hd__or2_1
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05765_ _11686_/Q _09998_/A _06924_/A _11733_/Q _06344_/C1 vssd1 vssd1 vccd1 vccd1
+ _05765_/X sky130_fd_sc_hd__o221a_1
X_08553_ _11129_/Q _08558_/S _07355_/S _07095_/B vssd1 vssd1 vccd1 vccd1 _11129_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07504_ _07796_/A _07504_/B vssd1 vssd1 vccd1 vccd1 _10536_/D sky130_fd_sc_hd__or2_1
XFILLER_51_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08484_ _09971_/A0 _08497_/S _08483_/X _08831_/C1 vssd1 vssd1 vccd1 vccd1 _11092_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05696_ _11109_/Q _05537_/Y _05573_/Y _11112_/Q _05695_/X vssd1 vssd1 vccd1 vccd1
+ _05704_/B sky130_fd_sc_hd__a221o_1
XFILLER_39_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07435_ _07143_/A _10494_/Q _07437_/S vssd1 vssd1 vccd1 vccd1 _07436_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07366_ _08733_/A _08051_/S vssd1 vssd1 vccd1 vccd1 _07373_/S sky130_fd_sc_hd__or2_4
XFILLER_109_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09105_ _11400_/Q _09243_/B _07591_/S _09192_/A vssd1 vssd1 vccd1 vccd1 _09105_/X
+ sky130_fd_sc_hd__a31o_1
X_06317_ _06287_/X _06900_/A _06299_/X _06316_/X vssd1 vssd1 vccd1 vccd1 _06317_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07297_ _07297_/A _07298_/B vssd1 vssd1 vccd1 vccd1 _07297_/Y sky130_fd_sc_hd__nor2_2
X_09036_ _10106_/A1 _09016_/X _09035_/X _09036_/C1 vssd1 vssd1 vccd1 vccd1 _11368_/D
+ sky130_fd_sc_hd__o211a_1
X_06248_ _11110_/Q _06737_/A2 _06736_/A2 _11196_/Q _06247_/X vssd1 vssd1 vccd1 vccd1
+ _06248_/X sky130_fd_sc_hd__o221a_1
XFILLER_136_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06179_ _11672_/Q _09391_/A _06284_/B1 _10997_/Q vssd1 vssd1 vccd1 vccd1 _06179_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout820 _09037_/A vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__buf_12
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout831 fanout846/X vssd1 vssd1 vccd1 vccd1 _06161_/A2 sky130_fd_sc_hd__buf_4
X_09938_ _11665_/Q _09938_/B vssd1 vssd1 vccd1 vccd1 _09938_/Y sky130_fd_sc_hd__nor2_1
Xfanout842 _09271_/A vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__buf_4
Xfanout853 fanout861/X vssd1 vssd1 vccd1 vccd1 _06371_/A2 sky130_fd_sc_hd__buf_4
Xfanout864 _05914_/A2 vssd1 vssd1 vccd1 vccd1 _07254_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_133_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout875 _10158_/A vssd1 vssd1 vccd1 vccd1 _06645_/A2 sky130_fd_sc_hd__clkbuf_16
Xfanout886 _06553_/B vssd1 vssd1 vccd1 vccd1 _06227_/A2 sky130_fd_sc_hd__buf_8
X_09869_ _09908_/A _09869_/B _09869_/C vssd1 vssd1 vccd1 vccd1 _09938_/B sky130_fd_sc_hd__or3_4
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout897 fanout901/X vssd1 vssd1 vccd1 vccd1 _06219_/A2 sky130_fd_sc_hd__clkbuf_8
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 _10021_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11762_/CLK _11762_/D vssd1 vssd1 vccd1 vccd1 _11762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10713_ _11458_/CLK _10713_/D vssd1 vssd1 vccd1 vccd1 _10713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11756_/CLK _11693_/D vssd1 vssd1 vccd1 vccd1 _11693_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10644_ _10644_/CLK _10644_/D vssd1 vssd1 vccd1 vccd1 _10644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10575_ _11458_/CLK _10575_/D vssd1 vssd1 vccd1 vccd1 _10575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127_ _11777_/CLK _11127_/D vssd1 vssd1 vccd1 vccd1 _11127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11058_ _11151_/CLK _11058_/D vssd1 vssd1 vccd1 vccd1 _11058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_wb_clk_i clkbuf_leaf_88_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11251_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10009_ _10009_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _10009_/Y sky130_fd_sc_hd__nor2_2
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05550_ _05616_/A1 _11429_/Q _11426_/Q _05077_/A vssd1 vssd1 vccd1 vccd1 _05550_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05481_ _10226_/Q input68/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05481_/X sky130_fd_sc_hd__mux2_1
X_07220_ _07039_/A _07776_/A2 _07771_/B1 _10377_/Q vssd1 vssd1 vccd1 vccd1 _10377_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07151_ _07151_/A _07151_/B _07151_/C _07151_/D vssd1 vssd1 vccd1 vccd1 _07151_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_9_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06102_ _11807_/Q _10180_/A _06100_/X _06101_/X vssd1 vssd1 vccd1 vccd1 _06102_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07082_ _07082_/A _08243_/C _08243_/D vssd1 vssd1 vccd1 vccd1 _08230_/B sky130_fd_sc_hd__or3_4
XFILLER_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06033_ _11512_/Q _09314_/A _06029_/X _06032_/X vssd1 vssd1 vccd1 vccd1 _06033_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_12_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07984_ _08196_/A _07984_/B vssd1 vssd1 vccd1 vccd1 _10816_/D sky130_fd_sc_hd__or2_1
XFILLER_86_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09723_ _11471_/Q _09883_/B1 _09953_/B1 _11477_/Q vssd1 vssd1 vccd1 vccd1 _09723_/X
+ sky130_fd_sc_hd__a22o_1
X_06935_ _10214_/Q _11568_/Q vssd1 vssd1 vccd1 vccd1 _06937_/B sky130_fd_sc_hd__xnor2_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09654_ _10354_/Q _09571_/B _09566_/C _10313_/Q _09653_/X vssd1 vssd1 vccd1 vccd1
+ _09659_/B sky130_fd_sc_hd__a221o_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06866_ _06861_/X _06862_/X _06865_/X _06860_/X vssd1 vssd1 vccd1 vccd1 _06866_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_82_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08605_ _10171_/A1 _11157_/Q _08621_/S vssd1 vssd1 vccd1 vccd1 _08606_/B sky130_fd_sc_hd__mux2_1
X_05817_ _05731_/X _06535_/A _05816_/X _06664_/C1 vssd1 vssd1 vccd1 vccd1 _05817_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06797_ _06853_/A1 _10245_/Q _06853_/A3 _06796_/X _05819_/B vssd1 vssd1 vccd1 vccd1
+ _06797_/X sky130_fd_sc_hd__a32o_1
X_09585_ _10507_/Q _09566_/A _09568_/D _10266_/Q _09580_/X vssd1 vssd1 vccd1 vccd1
+ _09586_/D sky130_fd_sc_hd__a221o_2
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05748_ _11867_/A _11868_/A _05751_/A vssd1 vssd1 vccd1 vccd1 _05748_/Y sky130_fd_sc_hd__nor3b_4
X_08536_ _08536_/A _08536_/B vssd1 vssd1 vccd1 vccd1 _11117_/D sky130_fd_sc_hd__or2_1
XFILLER_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08467_ _11085_/Q _08838_/A0 _08467_/S vssd1 vssd1 vccd1 vccd1 _08468_/B sky130_fd_sc_hd__mux2_1
X_05679_ _05679_/A _05679_/B _05679_/C _05679_/D vssd1 vssd1 vccd1 vccd1 _05680_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07418_ _07476_/A _07418_/B vssd1 vssd1 vccd1 vccd1 _10485_/D sky130_fd_sc_hd__or2_1
X_08398_ _11040_/Q _08422_/B vssd1 vssd1 vccd1 vccd1 _08398_/X sky130_fd_sc_hd__or2_1
XFILLER_143_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07349_ _10445_/Q _07350_/S _07846_/S _07333_/B vssd1 vssd1 vccd1 vccd1 _10445_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10360_ _11722_/CLK _10360_/D vssd1 vssd1 vccd1 vccd1 _10360_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09019_ _10182_/A0 _09035_/B _08664_/A vssd1 vssd1 vccd1 vccd1 _09019_/X sky130_fd_sc_hd__a21o_1
X_10291_ _11720_/CLK _10291_/D vssd1 vssd1 vccd1 vccd1 _10291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout650 _09497_/A vssd1 vssd1 vccd1 vccd1 _09492_/B sky130_fd_sc_hd__buf_4
Xfanout661 _11626_/Q vssd1 vssd1 vccd1 vccd1 _05077_/A sky130_fd_sc_hd__buf_8
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout672 _05349_/S vssd1 vssd1 vccd1 vccd1 _09680_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_150_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout683 _11598_/Q vssd1 vssd1 vccd1 vccd1 _05394_/S sky130_fd_sc_hd__buf_8
XFILLER_98_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout694 _05382_/S vssd1 vssd1 vccd1 vccd1 _05416_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11745_/CLK _11745_/D vssd1 vssd1 vccd1 vccd1 _11745_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11676_ _11685_/CLK _11676_/D vssd1 vssd1 vccd1 vccd1 _11676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10627_ _11474_/CLK _10627_/D vssd1 vssd1 vccd1 vccd1 _10627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10558_ _11575_/CLK _10558_/D vssd1 vssd1 vccd1 vccd1 _10558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10489_ _11711_/CLK _10489_/D vssd1 vssd1 vccd1 vccd1 _10489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06720_ _06720_/A _06720_/B vssd1 vssd1 vccd1 vccd1 _06720_/Y sky130_fd_sc_hd__nand2_2
X_06651_ _10369_/Q _09358_/A _09976_/A _10515_/Q _06651_/C1 vssd1 vssd1 vccd1 vccd1
+ _06651_/X sky130_fd_sc_hd__a221o_1
XFILLER_64_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05602_ _11682_/Q _05626_/A2 _05606_/B2 _11676_/Q _05601_/X vssd1 vssd1 vccd1 vccd1
+ _05603_/B sky130_fd_sc_hd__a221o_4
X_09370_ _10171_/A1 _09376_/B _10178_/B1 vssd1 vssd1 vccd1 vccd1 _09370_/X sky130_fd_sc_hd__a21o_1
X_06582_ _11283_/Q _09359_/A _09977_/A _10842_/Q _06624_/C1 vssd1 vssd1 vccd1 vccd1
+ _06582_/X sky130_fd_sc_hd__o221a_1
XFILLER_33_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05533_ _05629_/A2 _11526_/Q _11520_/Q _05629_/B1 vssd1 vssd1 vccd1 vccd1 _05533_/X
+ sky130_fd_sc_hd__a22o_1
X_08321_ _10118_/A0 _11000_/Q _08321_/S vssd1 vssd1 vccd1 vccd1 _11000_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08252_ _09985_/A1 _10958_/Q _08272_/S vssd1 vssd1 vccd1 vccd1 _08253_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05464_ _10755_/Q _09873_/B1 _09881_/B1 _10805_/Q _05461_/X vssd1 vssd1 vccd1 vccd1
+ _05466_/C sky130_fd_sc_hd__a221o_1
X_07203_ _07203_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _07205_/B sky130_fd_sc_hd__or2_4
X_08183_ _10925_/Q _07645_/B _07644_/Y _07229_/B vssd1 vssd1 vccd1 vccd1 _10925_/D
+ sky130_fd_sc_hd__o22a_1
X_05395_ _05395_/A _05395_/B _05395_/C _05395_/D vssd1 vssd1 vccd1 vccd1 _05401_/A
+ sky130_fd_sc_hd__or4_4
X_07134_ _07031_/A _07111_/X _07133_/X _07141_/B vssd1 vssd1 vccd1 vccd1 _10327_/D
+ sky130_fd_sc_hd__o211a_1
X_07065_ _10291_/Q _07078_/B vssd1 vssd1 vccd1 vccd1 _07065_/X sky130_fd_sc_hd__or2_1
X_06016_ _06450_/A _10225_/Q _06886_/A2 _06015_/X vssd1 vssd1 vccd1 vccd1 _10225_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07967_ _07441_/A _07966_/X _09241_/B1 vssd1 vssd1 vccd1 vccd1 _10806_/D sky130_fd_sc_hd__o21a_1
XFILLER_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09706_ _10416_/Q _09568_/A _09877_/B1 _10401_/Q _09705_/X vssd1 vssd1 vccd1 vccd1
+ _09713_/A sky130_fd_sc_hd__a221o_1
XFILLER_74_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06918_ _10200_/Q _06922_/B vssd1 vssd1 vccd1 vccd1 _06918_/X sky130_fd_sc_hd__or2_1
XFILLER_114_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07898_ _07147_/A _07966_/S _07897_/X _07902_/C1 vssd1 vssd1 vccd1 vccd1 _10767_/D
+ sky130_fd_sc_hd__o211a_1
X_09637_ _11658_/Q _11643_/Q vssd1 vssd1 vccd1 vccd1 _09637_/X sky130_fd_sc_hd__and2_1
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06849_ _10630_/Q _06860_/A2 _06848_/X _06849_/C1 vssd1 vssd1 vccd1 vccd1 _06849_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09568_ _09568_/A _09568_/B _09568_/C _09568_/D vssd1 vssd1 vccd1 vccd1 _09569_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_128_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08519_ _09285_/A1 _11109_/Q _08529_/S vssd1 vssd1 vccd1 vccd1 _08520_/B sky130_fd_sc_hd__mux2_1
XFILLER_145_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09499_ _09511_/C _09515_/B _09515_/C vssd1 vssd1 vccd1 vccd1 _09500_/C sky130_fd_sc_hd__and3b_1
XFILLER_19_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11530_ _11735_/CLK _11530_/D vssd1 vssd1 vccd1 vccd1 _11530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11461_ _11462_/CLK _11461_/D vssd1 vssd1 vccd1 vccd1 _11461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10412_ _11439_/CLK _10412_/D vssd1 vssd1 vccd1 vccd1 _10412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11392_ _11411_/CLK _11392_/D vssd1 vssd1 vccd1 vccd1 _11392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10343_ _11442_/CLK _10343_/D vssd1 vssd1 vccd1 vccd1 _10343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10274_ _11711_/CLK _10274_/D vssd1 vssd1 vccd1 vccd1 _10274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout480 _07205_/A vssd1 vssd1 vccd1 vccd1 _07147_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_63_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout491 _08843_/C1 vssd1 vssd1 vccd1 vccd1 _07003_/B sky130_fd_sc_hd__buf_4
XFILLER_47_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _11762_/CLK _11728_/D vssd1 vssd1 vccd1 vccd1 _11728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11659_ _11661_/CLK _11659_/D vssd1 vssd1 vccd1 vccd1 _11659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05180_ _10841_/Q _10840_/Q _05413_/S vssd1 vssd1 vccd1 vccd1 _05184_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08870_ _08987_/A1 _11292_/Q _08884_/S vssd1 vssd1 vccd1 vccd1 _08871_/B sky130_fd_sc_hd__mux2_1
XFILLER_97_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07821_ _07821_/A vssd1 vssd1 vccd1 vccd1 _07821_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07752_ _10677_/Q _07752_/B vssd1 vssd1 vccd1 vccd1 _07752_/X sky130_fd_sc_hd__or2_1
XFILLER_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06703_ _11617_/Q _06702_/X _06883_/B vssd1 vssd1 vccd1 vccd1 _10239_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07683_ _10639_/Q _07673_/Y _07676_/X _07016_/X vssd1 vssd1 vccd1 vccd1 _10639_/D
+ sky130_fd_sc_hd__a22o_1
X_09422_ _11652_/Q _11581_/Q _09704_/B vssd1 vssd1 vccd1 vccd1 _11581_/D sky130_fd_sc_hd__mux2_1
X_06634_ _10924_/Q _08166_/A _06634_/B1 _10446_/Q vssd1 vssd1 vccd1 vccd1 _06634_/X
+ sky130_fd_sc_hd__o22a_1
X_09353_ _10114_/A0 _11533_/Q _09357_/S vssd1 vssd1 vccd1 vccd1 _11533_/D sky130_fd_sc_hd__mux2_1
X_06565_ _10691_/Q _09358_/A _09976_/A _10514_/Q _07151_/A vssd1 vssd1 vccd1 vccd1
+ _06565_/X sky130_fd_sc_hd__a221o_1
XFILLER_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08304_ _08427_/A _08838_/S vssd1 vssd1 vccd1 vccd1 _08304_/Y sky130_fd_sc_hd__nand2_1
X_05516_ _05631_/A2 _10265_/Q _10261_/Q _05631_/B1 _05514_/X vssd1 vssd1 vccd1 vccd1
+ _05516_/X sky130_fd_sc_hd__a221o_1
X_09284_ _11494_/Q _09288_/B vssd1 vssd1 vccd1 vccd1 _09284_/X sky130_fd_sc_hd__or2_1
XFILLER_20_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06496_ _10830_/Q _07994_/A _06628_/B1 _11275_/Q vssd1 vssd1 vccd1 vccd1 _06496_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_60_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05447_ _10666_/Q _09568_/C _09573_/D _10659_/Q _05444_/X vssd1 vssd1 vccd1 vccd1
+ _05449_/C sky130_fd_sc_hd__a221o_1
X_08235_ _10951_/Q _08324_/B vssd1 vssd1 vccd1 vccd1 _08235_/X sky130_fd_sc_hd__or2_1
XFILLER_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08166_ _08166_/A _10119_/B _10119_/C vssd1 vssd1 vccd1 vccd1 _08166_/X sky130_fd_sc_hd__or3_4
X_05378_ _05378_/A _05378_/B _05378_/C _05378_/D vssd1 vssd1 vccd1 vccd1 _05379_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07117_ _10314_/Q _07126_/B _07123_/B1 _07229_/B vssd1 vssd1 vccd1 vccd1 _10314_/D
+ sky130_fd_sc_hd__o22a_1
X_08097_ _08097_/A _10119_/B _09038_/C vssd1 vssd1 vccd1 vccd1 _08097_/X sky130_fd_sc_hd__or3_2
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07048_ _07048_/A _10028_/A vssd1 vssd1 vccd1 vccd1 _07324_/B sky130_fd_sc_hd__and2_4
XFILLER_134_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08999_ _11351_/Q _09013_/B vssd1 vssd1 vccd1 vccd1 _08999_/X sky130_fd_sc_hd__or2_1
XFILLER_60_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_117_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11722_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10961_ _11319_/CLK _10961_/D vssd1 vssd1 vccd1 vccd1 _10961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10892_ _11601_/CLK _10892_/D vssd1 vssd1 vccd1 vccd1 _10892_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11513_ _11735_/CLK _11513_/D vssd1 vssd1 vccd1 vccd1 _11513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11444_ _11473_/CLK _11444_/D vssd1 vssd1 vccd1 vccd1 _11444_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_137_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11375_ _11410_/CLK _11375_/D vssd1 vssd1 vccd1 vccd1 _11375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10326_ _11745_/CLK _10326_/D vssd1 vssd1 vccd1 vccd1 _10326_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10257_ _11803_/CLK _10257_/D vssd1 vssd1 vccd1 vccd1 _10257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10188_ _07018_/A _11809_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _11809_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06350_ _10265_/Q _06976_/A _06903_/A _10202_/Q vssd1 vssd1 vccd1 vccd1 _06350_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05301_ _05301_/A _05301_/B _05301_/C _05301_/D vssd1 vssd1 vccd1 vccd1 _05302_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_148_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06281_ _11764_/Q _10108_/A _06279_/X _06280_/X vssd1 vssd1 vccd1 vccd1 _06281_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08020_ _10162_/A1 _08035_/S _08019_/X _07011_/B vssd1 vssd1 vccd1 vccd1 _10834_/D
+ sky130_fd_sc_hd__o211a_1
X_05232_ _05418_/S _10949_/Q vssd1 vssd1 vccd1 vccd1 _05232_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05163_ _11070_/Q _11069_/Q _05391_/S vssd1 vssd1 vccd1 vccd1 _05167_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09971_ _09971_/A0 _11671_/Q _09975_/S vssd1 vssd1 vccd1 vccd1 _11671_/D sky130_fd_sc_hd__mux2_1
X_05094_ _05819_/A vssd1 vssd1 vccd1 vccd1 _06892_/A sky130_fd_sc_hd__inv_12
XFILLER_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08922_ _11320_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08922_/X sky130_fd_sc_hd__or2_1
XFILLER_44_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08853_ _08853_/A1 _08850_/S _08852_/X _07011_/B vssd1 vssd1 vccd1 vccd1 _11284_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07804_ _07922_/A _07804_/B vssd1 vssd1 vccd1 vccd1 _10709_/D sky130_fd_sc_hd__or2_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08784_ _09101_/A1 _11248_/Q _08802_/S vssd1 vssd1 vccd1 vccd1 _08785_/B sky130_fd_sc_hd__mux2_1
X_05996_ _10438_/Q _06513_/A2 _06636_/A2 _11072_/Q _11869_/A vssd1 vssd1 vccd1 vccd1
+ _05996_/X sky130_fd_sc_hd__o221a_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07735_ _08939_/A1 _07761_/A2 _07734_/X _09201_/A1 vssd1 vssd1 vccd1 vccd1 _10668_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07666_ _10043_/A _07666_/B vssd1 vssd1 vccd1 vccd1 _10627_/D sky130_fd_sc_hd__or2_1
X_09405_ _11602_/Q _09554_/B vssd1 vssd1 vccd1 vccd1 _09406_/B sky130_fd_sc_hd__or2_4
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06617_ _11117_/Q _09081_/A _06613_/X _06616_/X vssd1 vssd1 vccd1 vccd1 _06617_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_0_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07597_ _07613_/A _08852_/B vssd1 vssd1 vccd1 vccd1 _07597_/Y sky130_fd_sc_hd__nor2_2
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09336_ _10168_/A1 _09326_/X _09335_/X _09993_/C1 vssd1 vssd1 vccd1 vccd1 _11522_/D
+ sky130_fd_sc_hd__o211a_1
X_06548_ _10449_/Q _07222_/A _07819_/A _10309_/Q vssd1 vssd1 vccd1 vccd1 _06552_/A
+ sky130_fd_sc_hd__o22a_1
X_09267_ _09995_/A1 _09249_/X _09266_/X _09267_/C1 vssd1 vssd1 vccd1 vccd1 _11486_/D
+ sky130_fd_sc_hd__o211a_1
X_06479_ _11467_/Q _06649_/A2 _06475_/X _06478_/X vssd1 vssd1 vccd1 vccd1 _06479_/X
+ sky130_fd_sc_hd__a211o_2
X_08218_ _08969_/A1 _08219_/S _08217_/X _08831_/C1 vssd1 vssd1 vccd1 vccd1 _10943_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09198_ _07243_/B _09193_/B _09191_/Y _11445_/Q _09193_/A vssd1 vssd1 vccd1 vccd1
+ _11445_/D sky130_fd_sc_hd__o221a_1
XFILLER_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08149_ _08469_/A _08140_/S _08148_/X _08345_/C1 vssd1 vssd1 vccd1 vccd1 _10900_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11160_ _11243_/CLK _11160_/D vssd1 vssd1 vccd1 vccd1 _11160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10111_ _10111_/A0 _11758_/Q _10118_/S vssd1 vssd1 vccd1 vccd1 _11758_/D sky130_fd_sc_hd__mux2_1
X_11091_ _11811_/CLK _11091_/D vssd1 vssd1 vccd1 vccd1 _11091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10042_ _11712_/Q _07028_/A _10057_/S vssd1 vssd1 vccd1 vccd1 _10043_/B sky130_fd_sc_hd__mux2_1
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10944_ _11312_/CLK _10944_/D vssd1 vssd1 vccd1 vccd1 _10944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10875_ _11777_/CLK _10875_/D vssd1 vssd1 vccd1 vccd1 _10875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_85_wb_clk_i clkbuf_leaf_85_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11330_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11776_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11427_ _11431_/CLK _11427_/D vssd1 vssd1 vccd1 vccd1 _11427_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_5 _05357_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ _11808_/CLK _11358_/D vssd1 vssd1 vccd1 vccd1 _11358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10309_ _11768_/CLK _10309_/D vssd1 vssd1 vccd1 vccd1 _10309_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11289_ _11325_/CLK _11289_/D vssd1 vssd1 vccd1 vccd1 _11289_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1050 _09280_/A1 vssd1 vssd1 vccd1 vccd1 _09141_/A1 sky130_fd_sc_hd__buf_6
Xfanout1061 _07785_/A0 vssd1 vssd1 vccd1 vccd1 _10166_/A1 sky130_fd_sc_hd__buf_8
XFILLER_120_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1072 input106/X vssd1 vssd1 vccd1 vccd1 _07036_/A sky130_fd_sc_hd__buf_6
X_05850_ _10747_/Q _07853_/A vssd1 vssd1 vccd1 vccd1 _05850_/X sky130_fd_sc_hd__or2_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05781_ _10554_/Q _07540_/A _06805_/B1 _10496_/Q vssd1 vssd1 vccd1 vccd1 _05781_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_47_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07520_ _07934_/A _07520_/B vssd1 vssd1 vccd1 vccd1 _10544_/D sky130_fd_sc_hd__or2_1
XFILLER_78_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07451_ _07451_/A _07451_/B vssd1 vssd1 vccd1 vccd1 _07451_/X sky130_fd_sc_hd__or2_4
XFILLER_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06402_ _11216_/Q _06126_/B _06398_/X _06401_/X vssd1 vssd1 vccd1 vccd1 _06402_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07382_ _10466_/Q _07015_/A _07393_/S vssd1 vssd1 vccd1 vccd1 _07383_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09121_ _11407_/Q _09127_/B vssd1 vssd1 vccd1 vccd1 _09121_/X sky130_fd_sc_hd__or2_1
X_06333_ _10738_/Q _06634_/B1 _06731_/B1 _11077_/Q _06550_/C1 vssd1 vssd1 vccd1 vccd1
+ _06333_/X sky130_fd_sc_hd__o221a_1
XFILLER_148_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09052_ _09285_/A1 _09038_/X _09051_/X _09289_/C1 vssd1 vssd1 vccd1 vccd1 _11375_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06264_ _10586_/Q _06454_/A2 _06455_/B1 _10430_/Q _06263_/X vssd1 vssd1 vccd1 vccd1
+ _06264_/X sky130_fd_sc_hd__o221a_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08003_ _09323_/A0 _10826_/Q _08011_/S vssd1 vssd1 vccd1 vccd1 _08004_/B sky130_fd_sc_hd__mux2_1
X_05215_ _10856_/Q _10855_/Q _05430_/S vssd1 vssd1 vccd1 vccd1 _05215_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_1284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06195_ _10687_/Q _07904_/A _06871_/A2 _10383_/Q vssd1 vssd1 vccd1 vccd1 _06195_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_116_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05146_ _05146_/A _05146_/B vssd1 vssd1 vccd1 vccd1 _05146_/Y sky130_fd_sc_hd__nor2_8
XFILLER_104_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05077_ _05077_/A vssd1 vssd1 vccd1 vccd1 _05077_/Y sky130_fd_sc_hd__clkinv_2
X_09954_ _10364_/Q _09566_/A _09568_/D _10682_/Q _09950_/X vssd1 vssd1 vccd1 vccd1
+ _09955_/D sky130_fd_sc_hd__a221o_1
XFILLER_89_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08905_ _07232_/B _08902_/C _08904_/X vssd1 vssd1 vccd1 vccd1 _11312_/D sky130_fd_sc_hd__a21o_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09885_ _11400_/Q _09568_/A _09565_/C _10568_/Q _09882_/X vssd1 vssd1 vccd1 vccd1
+ _09887_/C sky130_fd_sc_hd__a221o_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08836_ _11276_/Q _08840_/B vssd1 vssd1 vccd1 vccd1 _08836_/X sky130_fd_sc_hd__or2_1
XFILLER_131_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1104 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1104/HI io_oeb[34] sky130_fd_sc_hd__conb_1
X_08767_ _08869_/A _08767_/B vssd1 vssd1 vccd1 vccd1 _11239_/D sky130_fd_sc_hd__or2_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1115 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1115/HI io_out[7] sky130_fd_sc_hd__conb_1
X_05979_ _10381_/Q _06860_/A2 _06710_/B _10796_/Q vssd1 vssd1 vccd1 vccd1 _05979_/X
+ sky130_fd_sc_hd__o22a_1
Xwrapped_tms1x00_1126 vssd1 vssd1 vccd1 vccd1 io_oeb[3] wrapped_tms1x00_1126/LO sky130_fd_sc_hd__conb_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ _10660_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07718_/X sky130_fd_sc_hd__or2_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _08937_/A1 _08707_/S _08697_/X _08937_/C1 vssd1 vssd1 vccd1 vccd1 _11203_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07649_ _10613_/Q _07013_/X _07651_/S vssd1 vssd1 vccd1 vccd1 _10613_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ _11442_/CLK _10660_/D vssd1 vssd1 vccd1 vccd1 _10660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09319_ _10113_/A0 _11512_/Q _09324_/S vssd1 vssd1 vccd1 vccd1 _11512_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10591_ _11243_/CLK _10591_/D vssd1 vssd1 vccd1 vccd1 _10591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11212_ _11770_/CLK _11212_/D vssd1 vssd1 vccd1 vccd1 _11212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11143_ _11652_/CLK _11143_/D vssd1 vssd1 vccd1 vccd1 _11143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_132_wb_clk_i clkbuf_4_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11743_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11074_ _11177_/CLK _11074_/D vssd1 vssd1 vccd1 vccd1 _11074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10025_ _09214_/A _11703_/Q _10025_/S vssd1 vssd1 vccd1 vccd1 _10026_/B sky130_fd_sc_hd__mux2_1
XFILLER_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10927_ _10929_/CLK _10927_/D vssd1 vssd1 vccd1 vccd1 _10927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10858_ _11023_/CLK _10858_/D vssd1 vssd1 vccd1 vccd1 _10858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _11005_/CLK _10789_/D vssd1 vssd1 vccd1 vccd1 _10789_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout309 _07750_/B vssd1 vssd1 vccd1 vccd1 _07760_/B sky130_fd_sc_hd__buf_4
XFILLER_141_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06951_ _11662_/Q _05474_/B _06948_/X _05474_/A _06950_/X vssd1 vssd1 vccd1 vccd1
+ _06951_/X sky130_fd_sc_hd__a221o_4
XFILLER_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05902_ _11804_/Q _10180_/A _08097_/A _10195_/Q vssd1 vssd1 vccd1 vccd1 _05902_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09670_ _11633_/Q _09669_/Y _09447_/B vssd1 vssd1 vccd1 vccd1 _09670_/X sky130_fd_sc_hd__o21a_1
X_06882_ _10252_/Q _06883_/B _06883_/C vssd1 vssd1 vccd1 vccd1 _10252_/D sky130_fd_sc_hd__and3_1
XFILLER_67_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08621_ _08935_/A1 _11165_/Q _08621_/S vssd1 vssd1 vccd1 vccd1 _08622_/B sky130_fd_sc_hd__mux2_1
X_05833_ _11757_/Q _06161_/A2 _06284_/B1 _10992_/Q vssd1 vssd1 vccd1 vccd1 _05833_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_67_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08552_ _11128_/Q _08558_/S _07355_/S _07617_/B vssd1 vssd1 vccd1 vccd1 _11128_/D
+ sky130_fd_sc_hd__o22a_1
X_05764_ _11723_/Q _10061_/A _09347_/A _11528_/Q vssd1 vssd1 vccd1 vccd1 _05764_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07503_ _10021_/A0 _10536_/Q _07533_/S vssd1 vssd1 vccd1 vccd1 _07504_/B sky130_fd_sc_hd__mux2_1
XFILLER_63_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08483_ _11092_/Q _08503_/B vssd1 vssd1 vccd1 vccd1 _08483_/X sky130_fd_sc_hd__or2_1
XFILLER_23_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05695_ _11122_/Q _05518_/Y _05524_/Y _11113_/Q vssd1 vssd1 vccd1 vccd1 _05695_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07434_ _10058_/A _07434_/B vssd1 vssd1 vccd1 vccd1 _10493_/D sky130_fd_sc_hd__or2_1
XFILLER_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07365_ _08745_/A _08051_/S vssd1 vssd1 vccd1 vccd1 _07365_/Y sky130_fd_sc_hd__nor2_2
XFILLER_149_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09104_ _07451_/B _07539_/Y _09103_/X vssd1 vssd1 vccd1 vccd1 _11399_/D sky130_fd_sc_hd__a21o_1
XFILLER_109_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06316_ _06743_/B _06310_/X _06315_/X _07081_/A vssd1 vssd1 vccd1 vccd1 _06316_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07296_ _07039_/A _09187_/S _07295_/X _07902_/C1 vssd1 vssd1 vccd1 vccd1 _10416_/D
+ sky130_fd_sc_hd__o211a_1
X_09035_ _11368_/Q _09035_/B vssd1 vssd1 vccd1 vccd1 _09035_/X sky130_fd_sc_hd__or2_1
XFILLER_15_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06247_ _10962_/Q _06737_/B1 _08765_/A _11246_/Q vssd1 vssd1 vccd1 vccd1 _06247_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_102_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06178_ _11870_/A _06178_/B _06178_/C vssd1 vssd1 vccd1 vccd1 _06178_/X sky130_fd_sc_hd__or3_2
XFILLER_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05129_ _05129_/A _05129_/B _05129_/C _05129_/D vssd1 vssd1 vccd1 vccd1 _05135_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout810 _06766_/A2 vssd1 vssd1 vccd1 vccd1 _07152_/A sky130_fd_sc_hd__buf_8
XFILLER_85_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout821 _09037_/A vssd1 vssd1 vccd1 vccd1 _06649_/A2 sky130_fd_sc_hd__buf_12
XFILLER_137_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09937_ input9/X _09889_/Y _09926_/Y vssd1 vssd1 vccd1 vccd1 _09937_/X sky130_fd_sc_hd__a21o_1
Xfanout832 _06538_/A2 vssd1 vssd1 vccd1 vccd1 _06629_/A2 sky130_fd_sc_hd__buf_4
XFILLER_89_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout843 _06738_/A2 vssd1 vssd1 vccd1 vccd1 _09271_/A sky130_fd_sc_hd__buf_6
Xfanout854 _06459_/A2 vssd1 vssd1 vccd1 vccd1 _06630_/A2 sky130_fd_sc_hd__buf_4
Xfanout865 _05914_/A2 vssd1 vssd1 vccd1 vccd1 _06727_/B sky130_fd_sc_hd__buf_2
Xfanout876 _05740_/X vssd1 vssd1 vccd1 vccd1 _10158_/A sky130_fd_sc_hd__buf_12
XFILLER_133_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout887 fanout901/X vssd1 vssd1 vccd1 vccd1 _06553_/B sky130_fd_sc_hd__buf_8
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _09868_/A _09868_/B _09868_/C _09868_/D vssd1 vssd1 vccd1 vccd1 _09869_/C
+ sky130_fd_sc_hd__or4_2
Xfanout898 _06737_/A2 vssd1 vssd1 vccd1 vccd1 _09082_/A sky130_fd_sc_hd__buf_8
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08819_ _08819_/A _08819_/B vssd1 vssd1 vccd1 vccd1 _11267_/D sky130_fd_sc_hd__or2_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _10289_/Q _09947_/A2 _09947_/B1 _10294_/Q vssd1 vssd1 vccd1 vccd1 _09799_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _05401_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11765_/CLK _11761_/D vssd1 vssd1 vccd1 vccd1 _11761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10712_ _11458_/CLK _10712_/D vssd1 vssd1 vccd1 vccd1 _10712_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _11762_/CLK _11692_/D vssd1 vssd1 vccd1 vccd1 _11692_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10643_ _10644_/CLK _10643_/D vssd1 vssd1 vccd1 vccd1 _10643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10574_ _10782_/CLK _10574_/D vssd1 vssd1 vccd1 vccd1 _10574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11126_ _11268_/CLK _11126_/D vssd1 vssd1 vccd1 vccd1 _11126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11057_ _11269_/CLK _11057_/D vssd1 vssd1 vccd1 vccd1 _11057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10008_ _10118_/A0 _11695_/Q _10008_/S vssd1 vssd1 vccd1 vccd1 _11695_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05480_ _10225_/Q input67/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05480_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07150_ _10337_/Q _07150_/A2 _07188_/S _07043_/B vssd1 vssd1 vccd1 vccd1 _10337_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_125_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06101_ _10261_/Q _06976_/A _06903_/A _10198_/Q vssd1 vssd1 vccd1 vccd1 _06101_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07081_ _07081_/A _07151_/C _07151_/D vssd1 vssd1 vccd1 vccd1 _07643_/C sky130_fd_sc_hd__and3_4
XFILLER_12_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06032_ _11760_/Q _10108_/A _06030_/X _06031_/X vssd1 vssd1 vccd1 vccd1 _06032_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07983_ _10816_/Q _10128_/A0 _07991_/S vssd1 vssd1 vccd1 vccd1 _07984_/B sky130_fd_sc_hd__mux2_1
XFILLER_101_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09722_ _09908_/A _09722_/B vssd1 vssd1 vccd1 vccd1 _09722_/Y sky130_fd_sc_hd__nor2_2
X_06934_ _10106_/A1 _10212_/Q _06934_/S vssd1 vssd1 vccd1 vccd1 _10212_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09653_ _10311_/Q _09568_/D _09661_/B vssd1 vssd1 vccd1 vccd1 _09653_/X sky130_fd_sc_hd__a21bo_1
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06865_ _10416_/Q _07254_/A _06864_/X _06878_/C1 vssd1 vssd1 vccd1 vccd1 _06865_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08604_ _09141_/A1 _08621_/S _08603_/X _08791_/C1 vssd1 vssd1 vccd1 vccd1 _11156_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05816_ _05816_/A _05816_/B _05816_/C vssd1 vssd1 vccd1 vccd1 _05816_/X sky130_fd_sc_hd__or3_1
X_09584_ _10515_/Q _09944_/B1 _09948_/B1 _10272_/Q _09583_/X vssd1 vssd1 vccd1 vccd1
+ _09586_/C sky130_fd_sc_hd__a221o_2
X_06796_ _06853_/A1 _10245_/Q _06852_/A3 _06743_/X _06795_/X vssd1 vssd1 vccd1 vccd1
+ _06796_/X sky130_fd_sc_hd__a32o_1
XFILLER_55_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08535_ _09182_/A0 _11117_/Q _08537_/S vssd1 vssd1 vccd1 vccd1 _08536_/B sky130_fd_sc_hd__mux2_1
X_05747_ input79/X _11867_/A _11868_/A vssd1 vssd1 vccd1 vccd1 _05747_/Y sky130_fd_sc_hd__nand3_2
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08466_ _11084_/Q _08467_/S _08287_/Y _08817_/B2 vssd1 vssd1 vccd1 vccd1 _11084_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05678_ _11194_/Q _05609_/Y _05627_/Y _11189_/Q _05677_/X vssd1 vssd1 vccd1 vccd1
+ _05680_/C sky130_fd_sc_hd__a221o_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07417_ _07061_/A _10485_/Q _07429_/S vssd1 vssd1 vccd1 vccd1 _07418_/B sky130_fd_sc_hd__mux2_1
X_08397_ _08875_/A _08397_/B vssd1 vssd1 vccd1 vccd1 _11039_/D sky130_fd_sc_hd__or2_1
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07348_ _10444_/Q _07337_/X _07846_/S _07318_/B vssd1 vssd1 vccd1 vccd1 _10444_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07279_ _07028_/A _10408_/Q _09184_/S vssd1 vssd1 vccd1 vccd1 _07280_/B sky130_fd_sc_hd__mux2_1
XFILLER_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09018_ _10088_/A1 _09016_/X _09017_/X _09267_/C1 vssd1 vssd1 vccd1 vccd1 _11359_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10290_ _11706_/CLK _10290_/D vssd1 vssd1 vccd1 vccd1 _10290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout640 _05078_/Y vssd1 vssd1 vccd1 vccd1 _05630_/A2 sky130_fd_sc_hd__clkbuf_16
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout651 _09502_/A vssd1 vssd1 vccd1 vccd1 _09497_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout662 _11626_/Q vssd1 vssd1 vccd1 vccd1 _05628_/B1 sky130_fd_sc_hd__buf_6
XFILLER_120_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout673 _05349_/S vssd1 vssd1 vccd1 vccd1 _05397_/S sky130_fd_sc_hd__buf_8
XFILLER_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout684 _05300_/S vssd1 vssd1 vccd1 vccd1 _06945_/B sky130_fd_sc_hd__buf_8
XFILLER_150_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout695 _11596_/Q vssd1 vssd1 vccd1 vccd1 _05382_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11744_/CLK _11744_/D vssd1 vssd1 vccd1 vccd1 _11744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11675_ _11675_/CLK _11675_/D vssd1 vssd1 vccd1 vccd1 _11675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10626_ _11766_/CLK _10626_/D vssd1 vssd1 vccd1 vccd1 _10626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10557_ _11465_/CLK _10557_/D vssd1 vssd1 vccd1 vccd1 _10557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10488_ _11712_/CLK _10488_/D vssd1 vssd1 vccd1 vccd1 _10488_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11109_ _11319_/CLK _11109_/D vssd1 vssd1 vccd1 vccd1 _11109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06650_ _10291_/Q _09325_/A _09248_/A _10324_/Q vssd1 vssd1 vccd1 vccd1 _06650_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05601_ _11685_/Q _05631_/A2 _05631_/B1 _11681_/Q _05599_/X vssd1 vssd1 vccd1 vccd1
+ _05601_/X sky130_fd_sc_hd__a221o_1
XFILLER_91_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06581_ _10867_/Q _06976_/A _06903_/A _10907_/Q vssd1 vssd1 vccd1 vccd1 _06581_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_80_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08320_ _09323_/A0 _10999_/Q _08321_/S vssd1 vssd1 vccd1 vccd1 _10999_/D sky130_fd_sc_hd__mux2_1
X_05532_ _05628_/A2 _11525_/Q _11522_/Q _05628_/B1 vssd1 vssd1 vccd1 vccd1 _05532_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08251_ _08771_/A _08251_/B vssd1 vssd1 vccd1 vccd1 _10957_/D sky130_fd_sc_hd__or2_1
X_05463_ _10751_/Q _09877_/A2 _09886_/A2 _10749_/Q _05458_/X vssd1 vssd1 vccd1 vccd1
+ _05466_/B sky130_fd_sc_hd__a221o_1
X_07202_ _07202_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _07202_/Y sky130_fd_sc_hd__nor2_4
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08182_ _08647_/A _10924_/Q _08182_/S vssd1 vssd1 vccd1 vccd1 _10924_/D sky130_fd_sc_hd__mux2_1
X_05394_ _11216_/Q _11215_/Q _05394_/S vssd1 vssd1 vccd1 vccd1 _05395_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07133_ _10327_/Q _07145_/B vssd1 vssd1 vccd1 vccd1 _07133_/X sky130_fd_sc_hd__or2_1
X_07064_ _10050_/A _07064_/B vssd1 vssd1 vccd1 vccd1 _10290_/D sky130_fd_sc_hd__or2_1
XFILLER_134_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput210 _05485_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_4
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06015_ _05680_/X _06622_/A2 _06013_/X _06014_/Y vssd1 vssd1 vccd1 vccd1 _06015_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07966_ _08929_/A1 _10806_/Q _07966_/S vssd1 vssd1 vccd1 vccd1 _07966_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09705_ _10397_/Q _09875_/B1 _09886_/A2 _11433_/Q vssd1 vssd1 vccd1 vccd1 _09705_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06917_ _10150_/A1 _06903_/X _06916_/X _06990_/C1 vssd1 vssd1 vccd1 vccd1 _10199_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07897_ _10767_/Q _07901_/B vssd1 vssd1 vccd1 vccd1 _07897_/X sky130_fd_sc_hd__or2_1
XFILLER_114_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09636_ _09636_/A _09636_/B _09636_/C vssd1 vssd1 vccd1 vccd1 _09640_/B sky130_fd_sc_hd__or3_2
X_06848_ _10531_/Q _06873_/A2 _06871_/B1 _10736_/Q _06847_/X vssd1 vssd1 vccd1 vccd1
+ _06848_/X sky130_fd_sc_hd__o221a_1
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09567_ _09567_/A _09567_/B _09567_/C _09567_/D vssd1 vssd1 vccd1 vccd1 _09569_/C
+ sky130_fd_sc_hd__or4_1
X_06779_ _10714_/Q _07777_/A _07854_/A _10764_/Q _06778_/X vssd1 vssd1 vccd1 vccd1
+ _06779_/X sky130_fd_sc_hd__o221a_1
XFILLER_82_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08518_ _09283_/A1 _08529_/S _08517_/X _08919_/C1 vssd1 vssd1 vccd1 vccd1 _11108_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09498_ _11610_/Q _09496_/Y _09497_/X _09833_/A vssd1 vssd1 vccd1 vccd1 _11610_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08449_ _11070_/Q _07623_/X _07626_/S _07005_/A vssd1 vssd1 vccd1 vccd1 _11070_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_145_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11460_ _11474_/CLK _11460_/D vssd1 vssd1 vccd1 vccd1 _11460_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10411_ _10782_/CLK _10411_/D vssd1 vssd1 vccd1 vccd1 _10411_/Q sky130_fd_sc_hd__dfxtp_2
X_11391_ _11410_/CLK _11391_/D vssd1 vssd1 vccd1 vccd1 _11391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10342_ _11644_/CLK _10342_/D vssd1 vssd1 vccd1 vccd1 _10342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10273_ _11711_/CLK _10273_/D vssd1 vssd1 vccd1 vccd1 _10273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11763_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout470 _07018_/B vssd1 vssd1 vccd1 vccd1 _08662_/C1 sky130_fd_sc_hd__buf_6
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout481 fanout510/X vssd1 vssd1 vccd1 vccd1 _07205_/A sky130_fd_sc_hd__buf_8
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout492 _08843_/C1 vssd1 vssd1 vccd1 vccd1 _08791_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11762_/CLK _11727_/D vssd1 vssd1 vccd1 vccd1 _11727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11658_ _11661_/CLK _11658_/D vssd1 vssd1 vccd1 vccd1 _11658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10609_ _11777_/CLK _10609_/D vssd1 vssd1 vccd1 vccd1 _10609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11589_ _11650_/CLK _11589_/D vssd1 vssd1 vccd1 vccd1 _11589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07820_ _10039_/A _07820_/B vssd1 vssd1 vccd1 vccd1 _07820_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07751_ _07141_/A _07751_/A2 _07750_/X _07884_/C1 vssd1 vssd1 vccd1 vccd1 _10676_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06702_ _06695_/X _06700_/X _06701_/X vssd1 vssd1 vccd1 vccd1 _06702_/X sky130_fd_sc_hd__o21a_1
X_07682_ _10638_/Q _07674_/X _07675_/Y _07309_/X vssd1 vssd1 vccd1 vccd1 _10638_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09421_ _11651_/Q _11580_/Q _09704_/B vssd1 vssd1 vccd1 vccd1 _11580_/D sky130_fd_sc_hd__mux2_1
X_06633_ _06633_/A _06633_/B _06633_/C vssd1 vssd1 vccd1 vccd1 _06633_/X sky130_fd_sc_hd__or3_2
X_09352_ _10113_/A0 _11532_/Q _09357_/S vssd1 vssd1 vccd1 vccd1 _11532_/D sky130_fd_sc_hd__mux2_1
X_06564_ _10526_/Q _09325_/A _09248_/A _10322_/Q vssd1 vssd1 vccd1 vccd1 _06564_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08303_ _08303_/A _08840_/B vssd1 vssd1 vccd1 vccd1 _08303_/Y sky130_fd_sc_hd__nor2_1
X_05515_ _05630_/A2 _10259_/Q _10256_/Q _05079_/A _05513_/X vssd1 vssd1 vccd1 vccd1
+ _05518_/A sky130_fd_sc_hd__a221o_4
X_09283_ _09283_/A1 _09271_/X _09282_/X _09289_/C1 vssd1 vssd1 vccd1 vccd1 _11493_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06495_ _11611_/Q _06665_/A2 _06493_/B _06622_/B2 _06494_/X vssd1 vssd1 vccd1 vccd1
+ _10233_/D sky130_fd_sc_hd__a221o_1
XFILLER_127_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08234_ _09256_/A1 _08325_/B _08233_/X _08753_/C1 vssd1 vssd1 vccd1 vccd1 _10950_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05446_ _10660_/Q _09571_/B _09566_/C _10656_/Q _05438_/X vssd1 vssd1 vccd1 vccd1
+ _05449_/B sky130_fd_sc_hd__a221o_1
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08165_ _08853_/A1 _08162_/S _08164_/X _09993_/C1 vssd1 vssd1 vccd1 vccd1 _10908_/D
+ sky130_fd_sc_hd__o211a_1
X_05377_ _10827_/Q _10826_/Q _05377_/S vssd1 vssd1 vccd1 vccd1 _05378_/D sky130_fd_sc_hd__mux2_2
XFILLER_140_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07116_ _10313_/Q _07126_/B _07123_/B1 _07227_/B vssd1 vssd1 vccd1 vccd1 _10313_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08096_ _09292_/A _08649_/C _09037_/C vssd1 vssd1 vccd1 vccd1 _08362_/B sky130_fd_sc_hd__and3_4
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07047_ _07664_/A _07047_/B vssd1 vssd1 vccd1 vccd1 _07047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08998_ _10182_/A0 _08994_/X _08997_/X _09032_/C1 vssd1 vssd1 vccd1 vccd1 _11350_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07949_ _10791_/Q _07941_/Y _07944_/Y _09232_/B2 vssd1 vssd1 vccd1 vccd1 _10791_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10960_ _11291_/CLK _10960_/D vssd1 vssd1 vccd1 vccd1 _10960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09619_ _10737_/Q _09572_/A _09571_/D _10797_/Q vssd1 vssd1 vccd1 vccd1 _09626_/A
+ sky130_fd_sc_hd__a22o_1
X_10891_ _11604_/CLK _10891_/D vssd1 vssd1 vccd1 vccd1 _10891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11512_ _11735_/CLK _11512_/D vssd1 vssd1 vccd1 vccd1 _11512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11443_ _11450_/CLK _11443_/D vssd1 vssd1 vccd1 vccd1 _11443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11374_ _11410_/CLK _11374_/D vssd1 vssd1 vccd1 vccd1 _11374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10325_ _11719_/CLK _10325_/D vssd1 vssd1 vccd1 vccd1 _10325_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10256_ _11755_/CLK _10256_/D vssd1 vssd1 vccd1 vccd1 _10256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10187_ _08092_/A _11808_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _11808_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05300_ _11131_/Q _10447_/Q _05300_/S vssd1 vssd1 vccd1 vccd1 _05301_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06280_ _11731_/Q _10061_/A _09347_/A _11536_/Q vssd1 vssd1 vccd1 vccd1 _06280_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05231_ _05418_/S _11001_/Q vssd1 vssd1 vccd1 vccd1 _05231_/Y sky130_fd_sc_hd__nand2b_1
X_05162_ _05162_/A _05162_/B _05162_/C _05162_/D vssd1 vssd1 vccd1 vccd1 _05168_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09970_ _10113_/A0 _11670_/Q _09975_/S vssd1 vssd1 vccd1 vccd1 _11670_/D sky130_fd_sc_hd__mux2_1
X_05093_ input74/X vssd1 vssd1 vccd1 vccd1 _05093_/Y sky130_fd_sc_hd__inv_6
XFILLER_100_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08921_ _09285_/A1 _08945_/A2 _08920_/X _08921_/C1 vssd1 vssd1 vccd1 vccd1 _11319_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08852_ _11284_/Q _08852_/B vssd1 vssd1 vccd1 vccd1 _08852_/X sky130_fd_sc_hd__or2_1
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07803_ _08939_/A1 _10709_/Q _09193_/B vssd1 vssd1 vccd1 vccd1 _07804_/B sky130_fd_sc_hd__mux2_1
XFILLER_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08783_ _08783_/A _08783_/B vssd1 vssd1 vccd1 vccd1 _11247_/D sky130_fd_sc_hd__or2_1
X_05995_ _11126_/Q _06635_/A2 _08647_/B _11176_/Q vssd1 vssd1 vccd1 vccd1 _05995_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07734_ _10668_/Q _07760_/B vssd1 vssd1 vccd1 vccd1 _07734_/X sky130_fd_sc_hd__or2_1
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07665_ _10627_/Q _10047_/A1 _07665_/S vssd1 vssd1 vccd1 vccd1 _07666_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09404_ _11602_/Q _09554_/B vssd1 vssd1 vccd1 vccd1 _09404_/Y sky130_fd_sc_hd__nor2_4
X_06616_ _11166_/Q _09037_/A _06614_/X _06615_/X vssd1 vssd1 vccd1 vccd1 _06616_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07596_ _09359_/A _08665_/C _10159_/C vssd1 vssd1 vccd1 vccd1 _08850_/S sky130_fd_sc_hd__or3_4
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09335_ _11522_/Q _09343_/B vssd1 vssd1 vccd1 vccd1 _09335_/X sky130_fd_sc_hd__or2_1
X_06547_ _06538_/X _06539_/X _06541_/X _07689_/A vssd1 vssd1 vccd1 vccd1 _06547_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09266_ _11486_/Q _09266_/B vssd1 vssd1 vccd1 vccd1 _09266_/X sky130_fd_sc_hd__or2_1
XFILLER_90_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06478_ _10754_/Q _06648_/A2 _06477_/X _06873_/D1 vssd1 vssd1 vccd1 vccd1 _06478_/X
+ sky130_fd_sc_hd__a211o_1
X_08217_ _10943_/Q _08902_/C vssd1 vssd1 vccd1 vccd1 _08217_/X sky130_fd_sc_hd__or2_1
X_05429_ _11146_/Q _11145_/Q _05429_/S vssd1 vssd1 vccd1 vccd1 _05433_/A sky130_fd_sc_hd__mux2_1
X_09197_ _11444_/Q _09191_/Y _09192_/Y _07026_/X vssd1 vssd1 vccd1 vccd1 _11444_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08148_ _10900_/Q _08637_/C vssd1 vssd1 vccd1 vccd1 _08148_/X sky130_fd_sc_hd__or2_1
XFILLER_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08079_ _07059_/A _10865_/Q _08083_/S vssd1 vssd1 vccd1 vccd1 _08080_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10110_ _10110_/A0 _11757_/Q _10118_/S vssd1 vssd1 vccd1 vccd1 _11757_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11090_ _11607_/CLK _11090_/D vssd1 vssd1 vccd1 vccd1 _11090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10041_ _11711_/Q _10028_/B _10085_/S _07026_/B vssd1 vssd1 vccd1 vccd1 _11711_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10943_ _11312_/CLK _10943_/D vssd1 vssd1 vccd1 vccd1 _10943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10874_ _10939_/CLK _10874_/D vssd1 vssd1 vccd1 vccd1 _10874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11426_ _11801_/CLK _11426_/D vssd1 vssd1 vccd1 vccd1 _11426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _05379_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11005_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11357_ _11811_/CLK _11357_/D vssd1 vssd1 vccd1 vccd1 _11357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10308_ _10727_/CLK _10308_/D vssd1 vssd1 vccd1 vccd1 _10308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _11325_/CLK _11288_/D vssd1 vssd1 vccd1 vccd1 _11288_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _11663_/CLK _10239_/D vssd1 vssd1 vccd1 vccd1 _10239_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_121_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1040 _08919_/A1 vssd1 vssd1 vccd1 vccd1 _10149_/A1 sky130_fd_sc_hd__buf_8
Xfanout1051 _09280_/A1 vssd1 vssd1 vccd1 vccd1 _10168_/A1 sky130_fd_sc_hd__buf_4
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1062 input111/X vssd1 vssd1 vccd1 vccd1 _07785_/A0 sky130_fd_sc_hd__buf_6
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1073 input104/X vssd1 vssd1 vccd1 vccd1 _07076_/A sky130_fd_sc_hd__buf_8
XFILLER_86_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05780_ _10396_/Q _06804_/B _07455_/A _10654_/Q vssd1 vssd1 vccd1 vccd1 _05780_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_130_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07450_ _07036_/A _07535_/S _07442_/Y _10502_/Q _09193_/A vssd1 vssd1 vccd1 vccd1
+ _10502_/D sky130_fd_sc_hd__o221a_1
XFILLER_126_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06401_ _11264_/Q _06635_/B1 _06399_/X _06400_/X vssd1 vssd1 vccd1 vccd1 _06401_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07381_ _08733_/A _07381_/B vssd1 vssd1 vccd1 vccd1 _10465_/D sky130_fd_sc_hd__or2_1
XFILLER_76_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09120_ _11406_/Q _09110_/X _09119_/X vssd1 vssd1 vccd1 vccd1 _11406_/D sky130_fd_sc_hd__a21o_1
X_06332_ _10917_/Q _06591_/A2 _05865_/B _11774_/Q vssd1 vssd1 vccd1 vccd1 _06332_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09051_ _11375_/Q _09055_/B vssd1 vssd1 vccd1 vccd1 _09051_/X sky130_fd_sc_hd__or2_1
X_06263_ _11030_/Q _06413_/A2 _06539_/B1 _10837_/Q vssd1 vssd1 vccd1 vccd1 _06263_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08002_ _09971_/A0 _08015_/S _08001_/X _08831_/C1 vssd1 vssd1 vccd1 vccd1 _10825_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05214_ _05214_/A _05214_/B _05214_/C _05214_/D vssd1 vssd1 vccd1 vccd1 _05214_/Y
+ sky130_fd_sc_hd__nor4_4
XFILLER_129_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06194_ _10772_/Q _06194_/A2 _06193_/X _06651_/C1 vssd1 vssd1 vccd1 vccd1 _06194_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05145_ _05145_/A _05145_/B _05145_/C _05145_/D vssd1 vssd1 vccd1 vccd1 _05146_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05076_ _05076_/A vssd1 vssd1 vccd1 vccd1 _05076_/Y sky130_fd_sc_hd__inv_2
X_09953_ _10377_/Q _09568_/A _09953_/B1 _10378_/Q _09949_/X vssd1 vssd1 vccd1 vccd1
+ _09955_/C sky130_fd_sc_hd__a221o_2
XFILLER_98_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08904_ _11312_/Q _08323_/A _08219_/S _08303_/A vssd1 vssd1 vccd1 vccd1 _08904_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _10566_/Q _09884_/A2 _09567_/D _10569_/Q _09883_/X vssd1 vssd1 vccd1 vccd1
+ _09887_/B sky130_fd_sc_hd__a221o_1
XFILLER_44_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _08835_/A _08835_/B vssd1 vssd1 vccd1 vccd1 _11275_/D sky130_fd_sc_hd__or2_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _09111_/A1 _11239_/Q _08802_/S vssd1 vssd1 vccd1 vccd1 _08767_/B sky130_fd_sc_hd__mux2_1
Xwrapped_tms1x00_1105 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1105/HI io_oeb[35] sky130_fd_sc_hd__conb_1
X_05978_ _11433_/Q _06804_/B _06805_/B1 _10498_/Q _05975_/X vssd1 vssd1 vccd1 vccd1
+ _05978_/X sky130_fd_sc_hd__o221a_1
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapped_tms1x00_1116 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1116/HI io_out[8] sky130_fd_sc_hd__conb_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1127 vssd1 vssd1 vccd1 vccd1 io_oeb[4] wrapped_tms1x00_1127/LO sky130_fd_sc_hd__conb_1
X_07717_ _10021_/A0 _07751_/A2 _07716_/X _07894_/C1 vssd1 vssd1 vccd1 vccd1 _10659_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _11203_/Q _08705_/B vssd1 vssd1 vccd1 vccd1 _08697_/X sky130_fd_sc_hd__or2_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07648_ _10612_/Q _07008_/X _07651_/S vssd1 vssd1 vccd1 vccd1 _10612_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07579_ _08423_/A1 _10573_/Q _07593_/S vssd1 vssd1 vccd1 vccd1 _07580_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09318_ _10112_/A0 _11511_/Q _09324_/S vssd1 vssd1 vccd1 vccd1 _11511_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10590_ _11628_/CLK _10590_/D vssd1 vssd1 vccd1 vccd1 _10590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09249_ _09249_/A _09271_/B _10159_/C vssd1 vssd1 vccd1 vccd1 _09249_/X sky130_fd_sc_hd__or3_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11211_ _11770_/CLK _11211_/D vssd1 vssd1 vccd1 vccd1 _11211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11142_ _11629_/CLK _11142_/D vssd1 vssd1 vccd1 vccd1 _11142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11073_ _11177_/CLK _11073_/D vssd1 vssd1 vccd1 vccd1 _11073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput110 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 input110/X sky130_fd_sc_hd__buf_2
XFILLER_89_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10024_ _10026_/A _10024_/B vssd1 vssd1 vccd1 vccd1 _11702_/D sky130_fd_sc_hd__or2_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_101_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _10785_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10926_ _10929_/CLK _10926_/D vssd1 vssd1 vccd1 vccd1 _10926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10857_ _11601_/CLK _10857_/D vssd1 vssd1 vccd1 vccd1 _10857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _11234_/CLK _10788_/D vssd1 vssd1 vccd1 vccd1 _10788_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11409_ _11411_/CLK _11409_/D vssd1 vssd1 vccd1 vccd1 _11409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06950_ _06950_/A _06950_/B vssd1 vssd1 vccd1 vccd1 _06950_/X sky130_fd_sc_hd__and2_1
XFILLER_140_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05901_ _11758_/Q _10108_/A _05897_/X _05900_/X vssd1 vssd1 vccd1 vccd1 _05901_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06881_ _06883_/B _06881_/B vssd1 vssd1 vccd1 vccd1 _10251_/D sky130_fd_sc_hd__and2_1
X_08620_ _08847_/A _08620_/B vssd1 vssd1 vccd1 vccd1 _11164_/D sky130_fd_sc_hd__or2_1
X_05832_ _05824_/X _05826_/X _05831_/X vssd1 vssd1 vccd1 vccd1 _05832_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08551_ _11127_/Q _08558_/S _07355_/S _07229_/B vssd1 vssd1 vccd1 vccd1 _11127_/D
+ sky130_fd_sc_hd__o22a_1
X_05763_ _11666_/Q _09965_/A _08311_/A _10991_/Q vssd1 vssd1 vccd1 vccd1 _05763_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07502_ _07916_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _10535_/D sky130_fd_sc_hd__or2_1
XFILLER_51_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08482_ _08492_/A _08482_/B vssd1 vssd1 vccd1 vccd1 _11091_/D sky130_fd_sc_hd__or2_1
X_05694_ _11121_/Q _05591_/Y _05633_/Y _11104_/Q _05693_/X vssd1 vssd1 vccd1 vccd1
+ _05704_/A sky130_fd_sc_hd__a221o_1
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07433_ _07076_/A _10493_/Q _07437_/S vssd1 vssd1 vccd1 vccd1 _07434_/B sky130_fd_sc_hd__mux2_1
XFILLER_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07364_ _09325_/A _08649_/B _08560_/C vssd1 vssd1 vccd1 vccd1 _07364_/X sky130_fd_sc_hd__and3_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09103_ _11399_/Q _09243_/B _07591_/S _09192_/A vssd1 vssd1 vccd1 vccd1 _09103_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06315_ _11160_/Q _08594_/A _06311_/X _06314_/X vssd1 vssd1 vccd1 vccd1 _06315_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07295_ _10416_/Q _09175_/B vssd1 vssd1 vccd1 vccd1 _07295_/X sky130_fd_sc_hd__or2_1
X_09034_ _11367_/Q _09016_/X _09033_/X vssd1 vssd1 vccd1 vccd1 _11367_/D sky130_fd_sc_hd__a21o_1
X_06246_ _11320_/Q _06738_/A2 _06735_/B1 _11159_/Q vssd1 vssd1 vccd1 vccd1 _06246_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06177_ _11385_/Q _09060_/A _06173_/X _06176_/X vssd1 vssd1 vccd1 vccd1 _06178_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05128_ _10926_/Q _10925_/Q _05393_/S vssd1 vssd1 vccd1 vccd1 _05129_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout800 _06166_/A2 vssd1 vssd1 vccd1 vccd1 _06641_/A2 sky130_fd_sc_hd__buf_6
Xfanout811 _06166_/A2 vssd1 vssd1 vccd1 vccd1 _06766_/A2 sky130_fd_sc_hd__buf_6
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout822 _05744_/Y vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__buf_12
X_09936_ _11660_/Q _09770_/S _09934_/X _09935_/X vssd1 vssd1 vccd1 vccd1 _11660_/D
+ sky130_fd_sc_hd__o22a_1
Xfanout833 _05953_/A2 vssd1 vssd1 vccd1 vccd1 _06538_/A2 sky130_fd_sc_hd__buf_4
Xfanout844 _06413_/A2 vssd1 vssd1 vccd1 vccd1 _06738_/A2 sky130_fd_sc_hd__buf_6
XFILLER_86_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout855 _08200_/A vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__buf_6
Xfanout866 _05914_/A2 vssd1 vssd1 vccd1 vccd1 _06804_/B sky130_fd_sc_hd__buf_6
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout877 _06468_/B vssd1 vssd1 vccd1 vccd1 _06513_/A2 sky130_fd_sc_hd__buf_6
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _11448_/Q _09871_/A2 _09565_/D _10711_/Q _09866_/X vssd1 vssd1 vccd1 vccd1
+ _09868_/D sky130_fd_sc_hd__a221o_1
Xfanout888 _07904_/A vssd1 vssd1 vccd1 vccd1 _07203_/A sky130_fd_sc_hd__buf_6
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout899 _06737_/A2 vssd1 vssd1 vccd1 vccd1 _06716_/A2 sky130_fd_sc_hd__buf_4
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _11267_/Q _08818_/A1 _08820_/S vssd1 vssd1 vccd1 vccd1 _08819_/B sky130_fd_sc_hd__mux2_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09798_ _11652_/Q _08950_/B _09797_/X _09407_/A vssd1 vssd1 vccd1 vccd1 _11652_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_73_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _05401_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08749_ _08749_/A _08749_/B vssd1 vssd1 vccd1 vccd1 _11231_/D sky130_fd_sc_hd__or2_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11762_/CLK _11760_/D vssd1 vssd1 vccd1 vccd1 _11760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10711_ _10782_/CLK _10711_/D vssd1 vssd1 vccd1 vccd1 _10711_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11691_ _11765_/CLK _11691_/D vssd1 vssd1 vccd1 vccd1 _11691_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10642_ _11270_/CLK _10642_/D vssd1 vssd1 vccd1 vccd1 _10642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10573_ _10782_/CLK _10573_/D vssd1 vssd1 vccd1 vccd1 _10573_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11125_ _11177_/CLK _11125_/D vssd1 vssd1 vccd1 vccd1 _11125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11056_ _11269_/CLK _11056_/D vssd1 vssd1 vccd1 vccd1 _11056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10007_ _10117_/A0 _11694_/Q _10008_/S vssd1 vssd1 vccd1 vccd1 _11694_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10909_ _11766_/CLK _10909_/D vssd1 vssd1 vccd1 vccd1 _10909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06100_ _11364_/Q _09016_/A _08994_/A _11354_/Q _06349_/C1 vssd1 vssd1 vccd1 vccd1
+ _06100_/X sky130_fd_sc_hd__o221a_1
X_07080_ _10299_/Q _07078_/B _07496_/S _07040_/B vssd1 vssd1 vccd1 vccd1 _10299_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06031_ _11690_/Q _09998_/A _06924_/A _11737_/Q _06344_/C1 vssd1 vssd1 vccd1 vccd1
+ _06031_/X sky130_fd_sc_hd__o221a_1
XFILLER_114_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07982_ _10815_/Q _07977_/S _07363_/S _08811_/B2 vssd1 vssd1 vccd1 vccd1 _10815_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06933_ _10105_/A1 _10211_/Q _06934_/S vssd1 vssd1 vccd1 vccd1 _10211_/D sky130_fd_sc_hd__mux2_1
X_09721_ _09721_/A _09721_/B _09721_/C _09721_/D vssd1 vssd1 vccd1 vccd1 _09722_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_45_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06864_ _11449_/Q _07777_/A _07440_/A _10504_/Q _06863_/X vssd1 vssd1 vccd1 vccd1
+ _06864_/X sky130_fd_sc_hd__o221a_1
X_09652_ _10355_/Q _09571_/A _09572_/D _10317_/Q _09651_/X vssd1 vssd1 vccd1 vccd1
+ _09659_/A sky130_fd_sc_hd__a221o_1
XFILLER_55_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05815_ _07083_/A _05798_/X _05803_/X _05813_/X _06619_/A1 vssd1 vssd1 vccd1 vccd1
+ _05816_/C sky130_fd_sc_hd__o311a_1
XFILLER_94_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08603_ _11156_/Q _08633_/B vssd1 vssd1 vccd1 vccd1 _08603_/X sky130_fd_sc_hd__or2_1
X_09583_ _10517_/Q _09570_/A _09573_/C _10276_/Q vssd1 vssd1 vccd1 vccd1 _09583_/X
+ sky130_fd_sc_hd__a22o_1
X_06795_ _06790_/X _06791_/X _06794_/X _06789_/X vssd1 vssd1 vccd1 vccd1 _06795_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_24_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ _08793_/A _08534_/B vssd1 vssd1 vccd1 vccd1 _11116_/D sky130_fd_sc_hd__or2_1
X_05746_ _05751_/A _11867_/A _11868_/A vssd1 vssd1 vccd1 vccd1 _05746_/X sky130_fd_sc_hd__and3_4
X_08465_ _08749_/A _08465_/B vssd1 vssd1 vccd1 vccd1 _11083_/D sky130_fd_sc_hd__or2_1
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05677_ _11207_/Q _05591_/Y _05633_/Y _11190_/Q vssd1 vssd1 vccd1 vccd1 _05677_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07416_ _07420_/A _07416_/B vssd1 vssd1 vccd1 vccd1 _10484_/D sky130_fd_sc_hd__or2_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08396_ _09285_/A1 _11039_/Q _08404_/S vssd1 vssd1 vccd1 vccd1 _08397_/B sky130_fd_sc_hd__mux2_1
XFILLER_149_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07347_ _10443_/Q _07350_/S _07846_/S _07314_/B vssd1 vssd1 vccd1 vccd1 _10443_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07278_ _07796_/A _07278_/B vssd1 vssd1 vccd1 vccd1 _10407_/D sky130_fd_sc_hd__or2_1
XFILLER_136_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09017_ _11359_/Q _09035_/B vssd1 vssd1 vccd1 vccd1 _09017_/X sky130_fd_sc_hd__or2_1
X_06229_ _11366_/Q _10087_/A _08994_/A _11356_/Q _06349_/C1 vssd1 vssd1 vccd1 vccd1
+ _06229_/X sky130_fd_sc_hd__o221a_1
XFILLER_151_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout630 _05730_/Y vssd1 vssd1 vccd1 vccd1 _05819_/B sky130_fd_sc_hd__buf_12
XFILLER_28_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout641 _05078_/Y vssd1 vssd1 vccd1 vccd1 _05618_/A1 sky130_fd_sc_hd__buf_8
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09919_ _10477_/Q _09566_/C _09947_/B1 _10359_/Q _09918_/X vssd1 vssd1 vccd1 vccd1
+ _09919_/X sky130_fd_sc_hd__a221o_1
Xfanout652 _11656_/Q vssd1 vssd1 vccd1 vccd1 _09502_/A sky130_fd_sc_hd__buf_4
Xfanout663 _11625_/Q vssd1 vssd1 vccd1 vccd1 _05629_/B1 sky130_fd_sc_hd__buf_6
XFILLER_24_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout674 _06942_/B vssd1 vssd1 vccd1 vccd1 _05419_/S sky130_fd_sc_hd__buf_6
Xfanout685 _11598_/Q vssd1 vssd1 vccd1 vccd1 _05300_/S sky130_fd_sc_hd__buf_6
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout696 _05429_/S vssd1 vssd1 vccd1 vccd1 _05396_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _11812_/CLK _11812_/D vssd1 vssd1 vccd1 vccd1 _11812_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11743_/CLK _11743_/D vssd1 vssd1 vccd1 vccd1 _11743_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11674_ _11763_/CLK _11674_/D vssd1 vssd1 vccd1 vccd1 _11674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10625_ _10812_/CLK _10625_/D vssd1 vssd1 vccd1 vccd1 _10625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10556_ _11622_/CLK _10556_/D vssd1 vssd1 vccd1 vccd1 _10556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ _11712_/CLK _10487_/D vssd1 vssd1 vccd1 vccd1 _10487_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11108_ _11291_/CLK _11108_/D vssd1 vssd1 vccd1 vccd1 _11108_/Q sky130_fd_sc_hd__dfxtp_1
X_11039_ _11319_/CLK _11039_/D vssd1 vssd1 vccd1 vccd1 _11039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05600_ _11679_/Q _05630_/A2 _05620_/B2 _11677_/Q _05598_/X vssd1 vssd1 vccd1 vccd1
+ _05603_/A sky130_fd_sc_hd__a221o_4
X_06580_ _11237_/Q _07300_/A _09249_/A _11187_/Q vssd1 vssd1 vccd1 vccd1 _06580_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05531_ _05531_/A _05531_/B vssd1 vssd1 vccd1 vccd1 _05531_/Y sky130_fd_sc_hd__nor2_8
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08250_ _09364_/A1 _10957_/Q _08272_/S vssd1 vssd1 vccd1 vccd1 _08251_/B sky130_fd_sc_hd__mux2_1
XFILLER_75_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05462_ _10762_/Q _09879_/B1 _09948_/B1 _10756_/Q _05457_/X vssd1 vssd1 vccd1 vccd1
+ _05466_/A sky130_fd_sc_hd__a221o_2
XFILLER_20_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07201_ _07042_/A _07191_/B _07192_/A _10363_/Q _07451_/A vssd1 vssd1 vccd1 vccd1
+ _10363_/D sky130_fd_sc_hd__a221o_1
X_08181_ _08818_/A1 _10923_/Q _08181_/S vssd1 vssd1 vccd1 vccd1 _10923_/D sky130_fd_sc_hd__mux2_1
X_05393_ _11212_/Q _11211_/Q _05393_/S vssd1 vssd1 vccd1 vccd1 _05395_/C sky130_fd_sc_hd__mux2_1
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11651_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07132_ _10326_/Q _07150_/A2 _07188_/S _07241_/B vssd1 vssd1 vccd1 vccd1 _10326_/D
+ sky130_fd_sc_hd__o22a_1
X_07063_ _10134_/A0 _10290_/Q _07074_/S vssd1 vssd1 vccd1 vccd1 _07064_/B sky130_fd_sc_hd__mux2_1
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput200 _05505_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_4
Xoutput211 _05486_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_4
X_06014_ _05816_/A _05951_/Y _05820_/B vssd1 vssd1 vccd1 vccd1 _06014_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07965_ _07095_/B _07883_/B _07964_/X vssd1 vssd1 vccd1 vccd1 _10805_/D sky130_fd_sc_hd__a21o_1
X_09704_ _11602_/Q _09704_/B vssd1 vssd1 vccd1 vccd1 _09770_/S sky130_fd_sc_hd__nor2_8
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06916_ _10199_/Q _06922_/B vssd1 vssd1 vccd1 vccd1 _06916_/X sky130_fd_sc_hd__or2_1
XFILLER_96_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07896_ input106/X _07966_/S _07895_/X _07902_/C1 vssd1 vssd1 vccd1 vccd1 _10766_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09635_ _10726_/Q _09568_/C _09948_/B1 _10727_/Q _09634_/X vssd1 vssd1 vccd1 vccd1
+ _09636_/C sky130_fd_sc_hd__a221o_2
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06847_ _10335_/Q _06856_/A2 _06685_/B _11744_/Q vssd1 vssd1 vccd1 vccd1 _06847_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06778_ _10576_/Q _06877_/B1 _06875_/B1 _10675_/Q vssd1 vssd1 vccd1 vccd1 _06778_/X
+ sky130_fd_sc_hd__o22a_1
X_09566_ _09566_/A _09566_/B _09566_/C _09566_/D vssd1 vssd1 vccd1 vccd1 _09569_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08517_ _11108_/Q _08545_/B vssd1 vssd1 vccd1 vccd1 _08517_/X sky130_fd_sc_hd__or2_1
X_05729_ _05729_/A input87/X input78/X vssd1 vssd1 vccd1 vccd1 _05820_/B sky130_fd_sc_hd__and3_4
XFILLER_93_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09497_ _09497_/A _09502_/B _09495_/C vssd1 vssd1 vccd1 vccd1 _09497_/X sky130_fd_sc_hd__or3b_1
XFILLER_145_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08448_ _11069_/Q _08459_/S _07626_/S _07324_/B vssd1 vssd1 vccd1 vccd1 _11069_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ _08664_/A _08379_/B vssd1 vssd1 vccd1 vccd1 _11031_/D sky130_fd_sc_hd__or2_1
XFILLER_104_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ _10773_/CLK _10410_/D vssd1 vssd1 vccd1 vccd1 _10410_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11390_ _11393_/CLK _11390_/D vssd1 vssd1 vccd1 vccd1 _11390_/Q sky130_fd_sc_hd__dfxtp_1
X_10341_ _11465_/CLK _10341_/D vssd1 vssd1 vccd1 vccd1 _10341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10272_ _11710_/CLK _10272_/D vssd1 vssd1 vccd1 vccd1 _10272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout460 _07018_/B vssd1 vssd1 vccd1 vccd1 _08821_/A sky130_fd_sc_hd__buf_6
XFILLER_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout471 _10153_/C1 vssd1 vssd1 vccd1 vccd1 _09036_/C1 sky130_fd_sc_hd__buf_4
Xfanout482 _07882_/C1 vssd1 vssd1 vccd1 vccd1 _07902_/C1 sky130_fd_sc_hd__buf_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout493 fanout510/X vssd1 vssd1 vccd1 vccd1 _08843_/C1 sky130_fd_sc_hd__buf_4
XFILLER_150_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_79_wb_clk_i clkbuf_leaf_85_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11319_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11765_/CLK _11726_/D vssd1 vssd1 vccd1 vccd1 _11726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11657_ _11657_/CLK _11657_/D vssd1 vssd1 vccd1 vccd1 _11657_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10608_ _10932_/CLK _10608_/D vssd1 vssd1 vccd1 vccd1 _10608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11588_ _11650_/CLK _11588_/D vssd1 vssd1 vccd1 vccd1 _11588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10539_ _10804_/CLK _10539_/D vssd1 vssd1 vccd1 vccd1 _10539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07750_ _10676_/Q _07750_/B vssd1 vssd1 vccd1 vccd1 _07750_/X sky130_fd_sc_hd__or2_1
XFILLER_81_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06701_ _06577_/A _10239_/Q _06855_/B vssd1 vssd1 vccd1 vccd1 _06701_/X sky130_fd_sc_hd__a21o_1
XFILLER_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07681_ _10637_/Q _07673_/Y _07676_/X _07229_/X vssd1 vssd1 vccd1 vccd1 _10637_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09420_ _11650_/Q _11579_/Q _09704_/B vssd1 vssd1 vccd1 vccd1 _11579_/D sky130_fd_sc_hd__mux2_1
X_06632_ _10900_/Q _06632_/A2 _06628_/X _06631_/X vssd1 vssd1 vccd1 vccd1 _06633_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09351_ _10112_/A0 _11531_/Q _09357_/S vssd1 vssd1 vccd1 vccd1 _11531_/D sky130_fd_sc_hd__mux2_1
X_06563_ _10755_/Q _06648_/A2 _08971_/A _10567_/Q _06562_/X vssd1 vssd1 vccd1 vccd1
+ _06563_/X sky130_fd_sc_hd__a221o_4
XFILLER_80_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05514_ _05629_/A2 _10264_/Q _10258_/Q _05629_/B1 vssd1 vssd1 vccd1 vccd1 _05514_/X
+ sky130_fd_sc_hd__a22o_1
X_08302_ _08437_/A _08838_/S vssd1 vssd1 vccd1 vccd1 _08302_/Y sky130_fd_sc_hd__nand2_1
X_09282_ _11493_/Q _09288_/B vssd1 vssd1 vccd1 vccd1 _09282_/X sky130_fd_sc_hd__or2_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06494_ _06474_/X _06491_/X _06493_/X _06664_/C1 vssd1 vssd1 vccd1 vccd1 _06494_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08233_ _10950_/Q _08324_/B vssd1 vssd1 vccd1 vccd1 _08233_/X sky130_fd_sc_hd__or2_1
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05445_ _10673_/Q _09570_/A _09948_/B1 _10667_/Q _05439_/X vssd1 vssd1 vccd1 vccd1
+ _05449_/A sky130_fd_sc_hd__a221o_2
XFILLER_105_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08164_ _10908_/Q _08164_/B vssd1 vssd1 vccd1 vccd1 _08164_/X sky130_fd_sc_hd__or2_1
XFILLER_140_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05376_ _10833_/Q _10832_/Q _09680_/B vssd1 vssd1 vccd1 vccd1 _05378_/C sky130_fd_sc_hd__mux2_1
XFILLER_119_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07115_ _10312_/Q _07135_/A2 _07123_/B1 _07090_/A vssd1 vssd1 vccd1 vccd1 _10312_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_140_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08095_ _07232_/B _08091_/C _08094_/X vssd1 vssd1 vccd1 vccd1 _10872_/D sky130_fd_sc_hd__a21o_1
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07046_ _07046_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _07074_/S sky130_fd_sc_hd__or2_4
XFILLER_107_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08997_ _11350_/Q _09013_/B vssd1 vssd1 vccd1 vccd1 _08997_/X sky130_fd_sc_hd__or2_1
X_07948_ _10790_/Q _07941_/Y _07944_/Y _07016_/X vssd1 vssd1 vccd1 vccd1 _10790_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07879_ _10758_/Q _07893_/B vssd1 vssd1 vccd1 vccd1 _07879_/X sky130_fd_sc_hd__or2_1
XFILLER_141_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09618_ _09615_/X _09617_/X _09558_/A _09600_/Y vssd1 vssd1 vccd1 vccd1 _09618_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10890_ _11269_/CLK _10890_/D vssd1 vssd1 vccd1 vccd1 _10890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09549_ _11665_/Q _09538_/X _09542_/X vssd1 vssd1 vccd1 vccd1 _09549_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11511_ _11765_/CLK _11511_/D vssd1 vssd1 vccd1 vccd1 _11511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_126_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11702_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11442_ _11442_/CLK _11442_/D vssd1 vssd1 vccd1 vccd1 _11442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11373_ _11495_/CLK _11373_/D vssd1 vssd1 vccd1 vccd1 _11373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10324_ _11720_/CLK _10324_/D vssd1 vssd1 vccd1 vccd1 _10324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _10255_/CLK _10255_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10186_ _07052_/A _11807_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _11807_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout290 _08718_/S vssd1 vssd1 vccd1 vccd1 _08726_/S sky130_fd_sc_hd__buf_6
XFILLER_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11709_ _11716_/CLK _11709_/D vssd1 vssd1 vccd1 vccd1 _11709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05230_ _11004_/Q _10952_/Q _05414_/S vssd1 vssd1 vccd1 vccd1 _05230_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05161_ _11072_/Q _11071_/Q _05429_/S vssd1 vssd1 vccd1 vccd1 _05162_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05092_ _07690_/B vssd1 vssd1 vccd1 vccd1 _05092_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08920_ _11319_/Q _08946_/B vssd1 vssd1 vccd1 vccd1 _08920_/X sky130_fd_sc_hd__or2_1
XFILLER_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08851_ _08851_/A _08851_/B vssd1 vssd1 vccd1 vccd1 _11283_/D sky130_fd_sc_hd__or2_1
XFILLER_69_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07802_ _07922_/A _07802_/B vssd1 vssd1 vccd1 vccd1 _10708_/D sky130_fd_sc_hd__or2_1
XFILLER_84_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05994_ _11306_/Q _10010_/A _05990_/X _05993_/X vssd1 vssd1 vccd1 vccd1 _06000_/B
+ sky130_fd_sc_hd__o211a_1
X_08782_ _09172_/A1 _11247_/Q _08792_/S vssd1 vssd1 vccd1 vccd1 _08783_/B sky130_fd_sc_hd__mux2_1
X_07733_ _09182_/A0 _07761_/A2 _07732_/X _07932_/C1 vssd1 vssd1 vccd1 vccd1 _10667_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07664_ _07664_/A _07664_/B vssd1 vssd1 vccd1 vccd1 _10626_/D sky130_fd_sc_hd__or2_1
XFILLER_53_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09403_ _11603_/Q _11604_/Q vssd1 vssd1 vccd1 vccd1 _09403_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06615_ _11203_/Q _10158_/A _09292_/A _11253_/Q vssd1 vssd1 vccd1 vccd1 _06615_/X
+ sky130_fd_sc_hd__a22o_1
X_07595_ _09081_/A _08471_/B _10136_/C vssd1 vssd1 vccd1 vccd1 _08852_/B sky130_fd_sc_hd__and3_2
XFILLER_80_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09334_ _11521_/Q _09326_/X _09333_/X vssd1 vssd1 vccd1 vccd1 _11521_/D sky130_fd_sc_hd__a21o_1
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06546_ _10898_/Q _06632_/A2 _06542_/X _06545_/X vssd1 vssd1 vccd1 vccd1 _06546_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_55_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09265_ _10153_/A1 _09249_/X _09264_/X _09267_/C1 vssd1 vssd1 vccd1 vccd1 _11485_/D
+ sky130_fd_sc_hd__o211a_1
X_06477_ _10706_/Q _09059_/A _09109_/A _10540_/Q _06476_/X vssd1 vssd1 vccd1 vccd1
+ _06477_/X sky130_fd_sc_hd__a221o_2
X_05428_ _05428_/A _05428_/B _05428_/C _05428_/D vssd1 vssd1 vccd1 vccd1 _05434_/A
+ sky130_fd_sc_hd__or4_4
X_08216_ _10190_/A0 _08225_/S _08215_/X _08351_/C1 vssd1 vssd1 vccd1 vccd1 _10942_/D
+ sky130_fd_sc_hd__o211a_1
X_09196_ _11443_/Q _09191_/Y _09192_/Y _07105_/X vssd1 vssd1 vccd1 vccd1 _11443_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_140_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05359_ _10990_/Q _10989_/Q _05426_/S vssd1 vssd1 vccd1 vccd1 _05362_/B sky130_fd_sc_hd__mux2_1
X_08147_ _08839_/A _08147_/B vssd1 vssd1 vccd1 vccd1 _10899_/D sky130_fd_sc_hd__or2_1
XFILLER_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08078_ _10153_/A1 _08083_/S _08077_/X _08753_/C1 vssd1 vssd1 vccd1 vccd1 _10864_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07029_ _09214_/B _07241_/B vssd1 vssd1 vccd1 vccd1 _07029_/X sky130_fd_sc_hd__or2_1
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _11710_/Q _10028_/B _10085_/S _07211_/X vssd1 vssd1 vccd1 vccd1 _11710_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10942_ _11023_/CLK _10942_/D vssd1 vssd1 vccd1 vccd1 _10942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10873_ _11312_/CLK _10873_/D vssd1 vssd1 vccd1 vccd1 _10873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11425_ _11428_/CLK _11425_/D vssd1 vssd1 vccd1 vccd1 _11425_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_7 _05379_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11356_ _11366_/CLK _11356_/D vssd1 vssd1 vccd1 vccd1 _11356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10307_ _11777_/CLK _10307_/D vssd1 vssd1 vccd1 vccd1 _10307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11287_ _11385_/CLK _11287_/D vssd1 vssd1 vccd1 vccd1 _11287_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_94_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11473_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_156_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10238_ _11644_/CLK _10238_/D vssd1 vssd1 vccd1 vccd1 _10238_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1030 _08092_/A vssd1 vssd1 vccd1 vccd1 _10115_/A0 sky130_fd_sc_hd__buf_4
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1041 _08919_/A1 vssd1 vssd1 vccd1 vccd1 _07052_/A sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_23_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11151_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10169_ _11796_/Q _10159_/X _10168_/X vssd1 vssd1 vccd1 vccd1 _11796_/D sky130_fd_sc_hd__a21o_1
Xfanout1052 input112/X vssd1 vssd1 vccd1 vccd1 _09280_/A1 sky130_fd_sc_hd__buf_8
Xfanout1063 _08579_/A0 vssd1 vssd1 vccd1 vccd1 _10111_/A0 sky130_fd_sc_hd__buf_4
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1074 input103/X vssd1 vssd1 vccd1 vccd1 _07141_/A sky130_fd_sc_hd__buf_8
XFILLER_67_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06400_ _11131_/Q _07222_/A _07819_/A _10305_/Q vssd1 vssd1 vccd1 vccd1 _06400_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07380_ _10465_/Q _07052_/A _07380_/S vssd1 vssd1 vccd1 vccd1 _07381_/B sky130_fd_sc_hd__mux2_1
XFILLER_15_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06331_ _11225_/Q _08650_/A _06639_/B1 _10816_/Q _06330_/X vssd1 vssd1 vccd1 vccd1
+ _06331_/X sky130_fd_sc_hd__o221a_1
XFILLER_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09050_ _11374_/Q _09038_/X _09049_/X vssd1 vssd1 vccd1 vccd1 _11374_/D sky130_fd_sc_hd__a21o_1
X_06262_ _10422_/Q _06541_/A2 _06504_/B1 _11004_/Q vssd1 vssd1 vccd1 vccd1 _06262_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08001_ _10825_/Q _08091_/C vssd1 vssd1 vccd1 vccd1 _08001_/X sky130_fd_sc_hd__or2_1
X_05213_ _05213_/A _05213_/B _05213_/C _05213_/D vssd1 vssd1 vccd1 vccd1 _05214_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_141_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06193_ _10703_/Q _07778_/A _07853_/A _10805_/Q _06192_/X vssd1 vssd1 vccd1 vccd1
+ _06193_/X sky130_fd_sc_hd__o221a_2
XFILLER_11_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05144_ _10642_/Q _10641_/Q _06945_/B vssd1 vssd1 vccd1 vccd1 _05145_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05075_ _11628_/Q vssd1 vssd1 vccd1 vccd1 _05075_/Y sky130_fd_sc_hd__clkinv_2
X_09952_ _10685_/Q _09568_/B _09568_/C _10691_/Q _09945_/X vssd1 vssd1 vccd1 vccd1
+ _09955_/B sky130_fd_sc_hd__a221o_1
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08903_ _08092_/X _08219_/S _08902_/X _08427_/A vssd1 vssd1 vccd1 vccd1 _11311_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _10565_/Q _09573_/A _09883_/B1 _10572_/Q vssd1 vssd1 vccd1 vccd1 _09883_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08834_/A0 _11275_/Q _08838_/S vssd1 vssd1 vccd1 vccd1 _08835_/B sky130_fd_sc_hd__mux2_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08765_ _08765_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08765_/X sky130_fd_sc_hd__or2_4
X_05977_ _10700_/Q _07778_/A _07540_/A _10557_/Q _05974_/X vssd1 vssd1 vccd1 vccd1
+ _05977_/X sky130_fd_sc_hd__o221a_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_tms1x00_1106 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1106/HI io_oeb[36] sky130_fd_sc_hd__conb_1
XFILLER_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapped_tms1x00_1117 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1117/HI io_out[9] sky130_fd_sc_hd__conb_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1128 vssd1 vssd1 vccd1 vccd1 io_oeb[5] wrapped_tms1x00_1128/LO sky130_fd_sc_hd__conb_1
XFILLER_22_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07716_ _10659_/Q _07750_/B vssd1 vssd1 vccd1 vccd1 _07716_/X sky130_fd_sc_hd__or2_1
XFILLER_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08696_ _08773_/A _08696_/B vssd1 vssd1 vccd1 vccd1 _11202_/D sky130_fd_sc_hd__or2_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07647_ _10611_/Q _08326_/B2 _07651_/S vssd1 vssd1 vccd1 vccd1 _10611_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07578_ _07930_/A _07578_/B vssd1 vssd1 vccd1 vccd1 _10572_/D sky130_fd_sc_hd__or2_1
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09317_ _10111_/A0 _11510_/Q _09324_/S vssd1 vssd1 vccd1 vccd1 _11510_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06529_ _11325_/Q _06648_/A2 _09131_/A _11297_/Q _08243_/B vssd1 vssd1 vccd1 vccd1
+ _06529_/X sky130_fd_sc_hd__a221o_1
XFILLER_51_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09248_ _09248_/A _10158_/B _10158_/C vssd1 vssd1 vccd1 vccd1 _09266_/B sky130_fd_sc_hd__and3_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ _07614_/A _09187_/S _07232_/X vssd1 vssd1 vccd1 vccd1 _09179_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11210_ _11262_/CLK _11210_/D vssd1 vssd1 vccd1 vccd1 _11210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11141_ _11629_/CLK _11141_/D vssd1 vssd1 vccd1 vccd1 _11141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11072_ _11177_/CLK _11072_/D vssd1 vssd1 vccd1 vccd1 _11072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput100 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 input100/X sky130_fd_sc_hd__clkbuf_4
XFILLER_88_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput111 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 input111/X sky130_fd_sc_hd__clkbuf_8
XFILLER_62_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10023_ _10023_/A0 _11702_/Q _10025_/S vssd1 vssd1 vccd1 vccd1 _10024_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _10929_/CLK _10925_/D vssd1 vssd1 vccd1 vccd1 _10925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_141_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11268_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10856_ _10939_/CLK _10856_/D vssd1 vssd1 vccd1 vccd1 _10856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _11234_/CLK _10787_/D vssd1 vssd1 vccd1 vccd1 _10787_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11408_ _11411_/CLK _11408_/D vssd1 vssd1 vccd1 vccd1 _11408_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11339_ _11495_/CLK _11339_/D vssd1 vssd1 vccd1 vccd1 _11339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05900_ _11510_/Q _09314_/A _05898_/X _05899_/X vssd1 vssd1 vccd1 vccd1 _05900_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06880_ _10251_/Q _06883_/C _06879_/X _06743_/X vssd1 vssd1 vccd1 vccd1 _06881_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05831_ _05827_/X _05828_/X _05830_/X _07297_/A vssd1 vssd1 vccd1 vccd1 _05831_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05762_ _07297_/A _05762_/B _05762_/C vssd1 vssd1 vccd1 vccd1 _05762_/X sky130_fd_sc_hd__or3_2
X_08550_ _11126_/Q _08558_/S _07355_/S _07227_/B vssd1 vssd1 vccd1 vccd1 _11126_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07501_ _10019_/A0 _10535_/Q _07513_/S vssd1 vssd1 vccd1 vccd1 _07502_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05693_ _11108_/Q _05609_/Y _05627_/Y _11103_/Q vssd1 vssd1 vccd1 vccd1 _05693_/X
+ sky130_fd_sc_hd__a22o_1
X_08481_ _10113_/A0 _11091_/Q _08497_/S vssd1 vssd1 vccd1 vccd1 _08482_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07432_ _10058_/A _07432_/B vssd1 vssd1 vccd1 vccd1 _10492_/D sky130_fd_sc_hd__or2_1
XFILLER_50_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07363_ _08901_/A1 _10454_/Q _07363_/S vssd1 vssd1 vccd1 vccd1 _10454_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09102_ _11398_/Q _09082_/X _09101_/X vssd1 vssd1 vccd1 vccd1 _11398_/D sky130_fd_sc_hd__a21o_1
X_06314_ _11111_/Q _09082_/A _06312_/X _06313_/X vssd1 vssd1 vccd1 vccd1 _06314_/X
+ sky130_fd_sc_hd__o211a_1
X_07294_ _07147_/A _09187_/S _07293_/X _07882_/C1 vssd1 vssd1 vccd1 vccd1 _10415_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09033_ _10105_/A1 _09035_/B _08664_/A vssd1 vssd1 vccd1 vccd1 _09033_/X sky130_fd_sc_hd__a21o_1
X_06245_ _06240_/X _06241_/X _06244_/X _06239_/X vssd1 vssd1 vccd1 vccd1 _06245_/X
+ sky130_fd_sc_hd__a31o_1
X_06176_ _11428_/Q _08668_/A _06175_/X _06670_/D1 vssd1 vssd1 vccd1 vccd1 _06176_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05127_ _10613_/Q _10612_/Q _05396_/S vssd1 vssd1 vccd1 vccd1 _05129_/C sky130_fd_sc_hd__mux2_1
XFILLER_137_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout801 _06632_/A2 vssd1 vssd1 vccd1 vccd1 _08123_/A sky130_fd_sc_hd__buf_4
XFILLER_137_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09935_ _06962_/X _09908_/Y _09926_/Y vssd1 vssd1 vccd1 vccd1 _09935_/X sky130_fd_sc_hd__a21o_1
Xfanout812 _06412_/B1 vssd1 vssd1 vccd1 vccd1 _06539_/B1 sky130_fd_sc_hd__buf_4
Xfanout823 _06514_/A2 vssd1 vssd1 vccd1 vccd1 _06635_/B1 sky130_fd_sc_hd__buf_6
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout834 _05953_/A2 vssd1 vssd1 vccd1 vccd1 _10087_/A sky130_fd_sc_hd__clkbuf_8
Xfanout845 fanout846/X vssd1 vssd1 vccd1 vccd1 _06413_/A2 sky130_fd_sc_hd__buf_6
Xfanout856 _06459_/A2 vssd1 vssd1 vccd1 vccd1 _08200_/A sky130_fd_sc_hd__buf_4
Xfanout867 _06719_/A2 vssd1 vssd1 vccd1 vccd1 _05914_/A2 sky130_fd_sc_hd__buf_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _10700_/Q _09886_/A2 _09886_/B1 _11446_/Q vssd1 vssd1 vccd1 vccd1 _09866_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout878 _06553_/B vssd1 vssd1 vccd1 vccd1 _06468_/B sky130_fd_sc_hd__buf_6
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout889 _06194_/A2 vssd1 vssd1 vccd1 vccd1 _07904_/A sky130_fd_sc_hd__clkbuf_16
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08817_ _11266_/Q _08820_/S _07630_/Y _08817_/B2 vssd1 vssd1 vccd1 vccd1 _11266_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09797_ _11651_/Q _09404_/Y _09796_/X _09681_/B vssd1 vssd1 vccd1 vccd1 _09797_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _08838_/A0 _11231_/Q _08748_/S vssd1 vssd1 vccd1 vccd1 _08749_/B sky130_fd_sc_hd__mux2_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _10019_/A0 _11194_/Q _08695_/S vssd1 vssd1 vccd1 vccd1 _08680_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10710_ _11458_/CLK _10710_/D vssd1 vssd1 vccd1 vccd1 _10710_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11735_/CLK _11690_/D vssd1 vssd1 vccd1 vccd1 _11690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10641_ _10644_/CLK _10641_/D vssd1 vssd1 vccd1 vccd1 _10641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10572_ _10773_/CLK _10572_/D vssd1 vssd1 vccd1 vccd1 _10572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11124_ _11766_/CLK _11124_/D vssd1 vssd1 vccd1 vccd1 _11124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11055_ _11151_/CLK _11055_/D vssd1 vssd1 vccd1 vccd1 _11055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10006_ _10080_/A0 _11693_/Q _10008_/S vssd1 vssd1 vccd1 vccd1 _11693_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10908_ _11527_/CLK _10908_/D vssd1 vssd1 vccd1 vccd1 _10908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10839_ _11243_/CLK _10839_/D vssd1 vssd1 vccd1 vccd1 _10839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06030_ _11727_/Q _10061_/A _09347_/A _11532_/Q vssd1 vssd1 vccd1 vccd1 _06030_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07981_ _08733_/A _07981_/B vssd1 vssd1 vccd1 vccd1 _10814_/D sky130_fd_sc_hd__or2_1
XFILLER_113_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09720_ _11440_/Q _09953_/B1 _09565_/D _10410_/Q _09719_/X vssd1 vssd1 vccd1 vccd1
+ _09721_/D sky130_fd_sc_hd__a221o_1
X_06932_ _10153_/A1 _10210_/Q _06934_/S vssd1 vssd1 vccd1 vccd1 _10210_/D sky130_fd_sc_hd__mux2_1
XFILLER_45_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09651_ _10327_/Q _09567_/B _09565_/B _10321_/Q vssd1 vssd1 vccd1 vccd1 _09651_/X
+ sky130_fd_sc_hd__a22o_1
X_06863_ _11476_/Q _07153_/A _06877_/B1 _11400_/Q vssd1 vssd1 vccd1 vccd1 _06863_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08602_ _08847_/A _08602_/B vssd1 vssd1 vccd1 vccd1 _11155_/D sky130_fd_sc_hd__or2_1
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05814_ _05773_/X _05785_/X _05793_/X _07082_/A vssd1 vssd1 vccd1 vccd1 _05816_/B
+ sky130_fd_sc_hd__o31a_1
X_09582_ _10277_/Q _09567_/A _09566_/D _10522_/Q _09578_/X vssd1 vssd1 vccd1 vccd1
+ _09586_/B sky130_fd_sc_hd__a221o_2
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06794_ _10785_/Q _06862_/A2 _06793_/X _06808_/C1 vssd1 vssd1 vccd1 vccd1 _06794_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08533_ _08883_/A1 _11116_/Q _08537_/S vssd1 vssd1 vccd1 vccd1 _08534_/B sky130_fd_sc_hd__mux2_1
X_05745_ _05745_/A _05749_/A _05751_/B vssd1 vssd1 vccd1 vccd1 _05745_/X sky130_fd_sc_hd__or3b_4
XFILLER_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08464_ _11083_/Q _08834_/A0 _08467_/S vssd1 vssd1 vccd1 vccd1 _08465_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_05676_ _11192_/Q _05567_/Y _05621_/Y _11201_/Q vssd1 vssd1 vccd1 vccd1 _05679_/D
+ sky130_fd_sc_hd__a22o_1
X_07415_ _07059_/A _10484_/Q _07429_/S vssd1 vssd1 vccd1 vccd1 _07416_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08395_ _08869_/A _08395_/B vssd1 vssd1 vccd1 vccd1 _11038_/D sky130_fd_sc_hd__or2_1
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ _10442_/Q _07350_/S _07346_/B1 _08811_/B2 vssd1 vssd1 vccd1 vccd1 _10442_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07277_ _09216_/A0 _10407_/Q _07277_/S vssd1 vssd1 vccd1 vccd1 _07278_/B sky130_fd_sc_hd__mux2_1
XFILLER_104_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09016_ _09016_/A _10180_/C _10137_/B vssd1 vssd1 vccd1 vccd1 _09016_/X sky130_fd_sc_hd__or3_4
X_06228_ _11565_/Q _06228_/A2 _09380_/A _11555_/Q vssd1 vssd1 vccd1 vccd1 _06228_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06159_ _11059_/Q _08054_/A _08123_/A _11173_/Q _06392_/C1 vssd1 vssd1 vccd1 vccd1
+ _06159_/X sky130_fd_sc_hd__o221a_1
XFILLER_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout620 _06748_/A2 vssd1 vssd1 vccd1 vccd1 _06807_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout631 _09478_/A vssd1 vssd1 vccd1 vccd1 _09407_/A sky130_fd_sc_hd__buf_6
Xfanout642 _05619_/B2 vssd1 vssd1 vccd1 vccd1 _05631_/B1 sky130_fd_sc_hd__buf_6
X_09918_ _10475_/Q _09568_/D _09948_/B1 _10486_/Q vssd1 vssd1 vccd1 vccd1 _09918_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout653 _09511_/C vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__clkbuf_4
Xfanout664 _11625_/Q vssd1 vssd1 vccd1 vccd1 _05078_/A sky130_fd_sc_hd__buf_8
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout675 _05349_/S vssd1 vssd1 vccd1 vccd1 _06942_/B sky130_fd_sc_hd__buf_6
Xfanout686 _05326_/S vssd1 vssd1 vccd1 vccd1 _05426_/S sky130_fd_sc_hd__buf_8
X_09849_ _11462_/Q _09568_/A _09565_/D _10782_/Q _09848_/X vssd1 vssd1 vccd1 vccd1
+ _09850_/D sky130_fd_sc_hd__a221o_1
XFILLER_24_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout697 _11595_/Q vssd1 vssd1 vccd1 vccd1 _05429_/S sky130_fd_sc_hd__buf_12
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11811_/CLK _11811_/D vssd1 vssd1 vccd1 vccd1 _11811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11742_ _11765_/CLK _11742_/D vssd1 vssd1 vccd1 vccd1 _11742_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11735_/CLK _11673_/D vssd1 vssd1 vccd1 vccd1 _11673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10624_ _10727_/CLK _10624_/D vssd1 vssd1 vccd1 vccd1 _10624_/Q sky130_fd_sc_hd__dfxtp_1
X_10555_ _11622_/CLK _10555_/D vssd1 vssd1 vccd1 vccd1 _10555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10486_ _11710_/CLK _10486_/D vssd1 vssd1 vccd1 vccd1 _10486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11107_ _11330_/CLK _11107_/D vssd1 vssd1 vccd1 vccd1 _11107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11038_ _11291_/CLK _11038_/D vssd1 vssd1 vccd1 vccd1 _11038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05530_ _05626_/A2 _11504_/Q _11499_/Q _05630_/B1 _05529_/X vssd1 vssd1 vccd1 vccd1
+ _05531_/B sky130_fd_sc_hd__a221o_4
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05461_ _10765_/Q _09876_/A2 _09874_/A2 _10746_/Q vssd1 vssd1 vccd1 vccd1 _05461_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07200_ _07039_/A _07191_/B _07192_/A _10362_/Q _07451_/A vssd1 vssd1 vccd1 vccd1
+ _10362_/D sky130_fd_sc_hd__a221o_1
XFILLER_60_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05392_ _11214_/Q _11213_/Q _05392_/S vssd1 vssd1 vccd1 vccd1 _05395_/B sky130_fd_sc_hd__mux2_1
X_08180_ _08661_/A _10922_/Q _08181_/S vssd1 vssd1 vccd1 vccd1 _10922_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07131_ _07025_/A _07111_/X _07130_/X _07147_/B vssd1 vssd1 vccd1 vccd1 _10325_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07062_ _10289_/Q _07047_/B _07490_/S _07318_/B vssd1 vssd1 vccd1 vccd1 _10289_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput201 _05506_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_4
X_06013_ _05787_/X _06011_/X _06012_/X _05816_/A vssd1 vssd1 vccd1 vccd1 _06013_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_138_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07964_ _10805_/Q _09206_/A _07871_/S _07599_/A vssd1 vssd1 vccd1 vccd1 _07964_/X
+ sky130_fd_sc_hd__a31o_1
X_09703_ _09703_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _11642_/D sky130_fd_sc_hd__or2_1
XFILLER_101_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06915_ _10198_/Q _06903_/X _06914_/X vssd1 vssd1 vccd1 vccd1 _10198_/D sky130_fd_sc_hd__a21o_1
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07895_ _10766_/Q _07901_/B vssd1 vssd1 vccd1 vccd1 _07895_/X sky130_fd_sc_hd__or2_1
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09634_ _10728_/Q _09944_/B1 _09947_/B1 _10800_/Q _09620_/X vssd1 vssd1 vccd1 vccd1
+ _09634_/X sky130_fd_sc_hd__a221o_1
XFILLER_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06846_ _10376_/Q _07904_/A _06870_/B1 _10522_/Q vssd1 vssd1 vccd1 vccd1 _06846_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09565_ _09565_/A _09565_/B _09565_/C _09565_/D vssd1 vssd1 vccd1 vccd1 _09569_/A
+ sky130_fd_sc_hd__or4_1
X_06777_ _10352_/Q _07153_/A _07440_/A _10549_/Q vssd1 vssd1 vccd1 vccd1 _06777_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08516_ _09280_/A1 _08537_/S _08515_/X _07003_/B vssd1 vssd1 vccd1 vccd1 _11107_/D
+ sky130_fd_sc_hd__o211a_1
X_05728_ _05728_/A _05728_/B _05728_/C _05728_/D vssd1 vssd1 vccd1 vccd1 _05728_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_145_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09496_ _09496_/A vssd1 vssd1 vccd1 vccd1 _09496_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08447_ _11068_/Q _08437_/Y _08438_/Y _07335_/X vssd1 vssd1 vccd1 vccd1 _11068_/D
+ sky130_fd_sc_hd__o22a_1
X_05659_ _11242_/Q _05567_/Y _05621_/Y _11251_/Q vssd1 vssd1 vccd1 vccd1 _05661_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08378_ _08760_/A0 _11031_/Q _08439_/B vssd1 vssd1 vccd1 vccd1 _08379_/B sky130_fd_sc_hd__mux2_1
XFILLER_149_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07329_ _10429_/Q _07322_/Y _07326_/Y _07229_/X vssd1 vssd1 vccd1 vccd1 _10429_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10340_ _11442_/CLK _10340_/D vssd1 vssd1 vccd1 vccd1 _10340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10271_ _11702_/CLK _10271_/D vssd1 vssd1 vccd1 vccd1 _10271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout450 _05146_/Y vssd1 vssd1 vccd1 vccd1 _09571_/B sky130_fd_sc_hd__buf_6
Xfanout461 _07107_/B vssd1 vssd1 vccd1 vccd1 _10028_/A sky130_fd_sc_hd__buf_8
XFILLER_63_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout472 _10153_/C1 vssd1 vssd1 vccd1 vccd1 _09032_/C1 sky130_fd_sc_hd__buf_2
XFILLER_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout483 _09201_/A1 vssd1 vssd1 vccd1 vccd1 _07932_/C1 sky130_fd_sc_hd__buf_4
Xfanout494 _09993_/C1 vssd1 vssd1 vccd1 vccd1 _09995_/C1 sky130_fd_sc_hd__buf_4
XFILLER_24_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _11735_/CLK _11725_/D vssd1 vssd1 vccd1 vccd1 _11725_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_48_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11485_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11656_ _11663_/CLK _11656_/D vssd1 vssd1 vccd1 vccd1 _11656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10607_ _10932_/CLK _10607_/D vssd1 vssd1 vccd1 vccd1 _10607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11587_ _11634_/CLK _11587_/D vssd1 vssd1 vccd1 vccd1 _11587_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10538_ _10666_/CLK _10538_/D vssd1 vssd1 vccd1 vccd1 _10538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10469_ _11629_/CLK _10469_/D vssd1 vssd1 vccd1 vccd1 _10469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06700_ _06696_/X _06697_/X _06699_/X _06852_/A3 vssd1 vssd1 vccd1 vccd1 _06700_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_38_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07680_ _10636_/Q _07673_/Y _07676_/X _07227_/X vssd1 vssd1 vccd1 vccd1 _10636_/D
+ sky130_fd_sc_hd__a22o_1
X_06631_ _10860_/Q _06631_/A2 _06629_/X _06630_/X vssd1 vssd1 vccd1 vccd1 _06631_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09350_ _10111_/A0 _11530_/Q _09357_/S vssd1 vssd1 vccd1 vccd1 _11530_/D sky130_fd_sc_hd__mux2_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06562_ _10707_/Q _09059_/A _09131_/A _10666_/Q _06561_/X vssd1 vssd1 vccd1 vccd1
+ _06562_/X sky130_fd_sc_hd__a221o_1
X_08301_ _08655_/B _08840_/B vssd1 vssd1 vccd1 vccd1 _08301_/Y sky130_fd_sc_hd__nor2_1
X_05513_ _05628_/A2 _10263_/Q _10260_/Q _05628_/B1 vssd1 vssd1 vccd1 vccd1 _05513_/X
+ sky130_fd_sc_hd__a22o_1
X_09281_ _11492_/Q _09271_/X _09280_/X vssd1 vssd1 vccd1 vccd1 _11492_/D sky130_fd_sc_hd__a21o_1
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06493_ _06855_/B _06493_/B vssd1 vssd1 vccd1 vccd1 _06493_/X sky130_fd_sc_hd__or2_1
XFILLER_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08232_ _10088_/A1 _08325_/B _08231_/X _08753_/C1 vssd1 vssd1 vccd1 vccd1 _10949_/D
+ sky130_fd_sc_hd__o211a_1
X_05444_ _10677_/Q _09571_/A _09566_/A _10654_/Q vssd1 vssd1 vccd1 vccd1 _05444_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08163_ _08761_/A _08163_/B vssd1 vssd1 vccd1 vccd1 _10907_/D sky130_fd_sc_hd__or2_1
X_05375_ _10831_/Q _10830_/Q _09680_/C vssd1 vssd1 vccd1 vccd1 _05378_/B sky130_fd_sc_hd__mux2_2
XFILLER_147_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07114_ _10311_/Q _07135_/A2 _07186_/S _07225_/A vssd1 vssd1 vccd1 vccd1 _10311_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_88_1336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ _10872_/Q _08437_/A _08011_/S _08303_/A vssd1 vssd1 vccd1 vccd1 _08094_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07045_ _07046_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _07045_/Y sky130_fd_sc_hd__nor2_4
XFILLER_133_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08996_ _10088_/A1 _08994_/X _08995_/X _09267_/C1 vssd1 vssd1 vccd1 vccd1 _11349_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07947_ _10789_/Q _07941_/Y _07944_/Y _07617_/X vssd1 vssd1 vccd1 vccd1 _10789_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07878_ _08939_/A1 _07871_/S _07877_/X _07884_/C1 vssd1 vssd1 vccd1 vccd1 _10757_/D
+ sky130_fd_sc_hd__o211a_1
X_09617_ _09617_/A _09617_/B _09617_/C _09617_/D vssd1 vssd1 vccd1 vccd1 _09617_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06829_ _10298_/Q _06873_/A2 _06710_/B _10802_/Q _06828_/X vssd1 vssd1 vccd1 vccd1
+ _06829_/X sky130_fd_sc_hd__o221a_1
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09548_ _05077_/A _09541_/Y _09547_/X _09833_/A vssd1 vssd1 vccd1 vccd1 _11626_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09479_ _11602_/Q _08950_/B _11603_/Q vssd1 vssd1 vccd1 vccd1 _09479_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _11735_/CLK _11510_/D vssd1 vssd1 vccd1 vccd1 _11510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11441_ _11442_/CLK _11441_/D vssd1 vssd1 vccd1 vccd1 _11441_/Q sky130_fd_sc_hd__dfxtp_1
X_11372_ _11410_/CLK _11372_/D vssd1 vssd1 vccd1 vccd1 _11372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10323_ _11706_/CLK _10323_/D vssd1 vssd1 vccd1 vccd1 _10323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10254_ _10255_/CLK hold1/X vssd1 vssd1 vccd1 vccd1 _10254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10185_ _10185_/A0 _11806_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _11806_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout280 _09206_/B vssd1 vssd1 vccd1 vccd1 _09221_/C sky130_fd_sc_hd__buf_8
Xfanout291 _07839_/A2 vssd1 vssd1 vccd1 vccd1 _07820_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11716_/CLK _11708_/D vssd1 vssd1 vccd1 vccd1 _11708_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11639_ _11652_/CLK _11639_/D vssd1 vssd1 vccd1 vccd1 _11639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05160_ _10599_/Q _11079_/Q _05397_/S vssd1 vssd1 vccd1 vccd1 _05162_/C sky130_fd_sc_hd__mux2_1
XFILLER_155_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05091_ _11870_/A vssd1 vssd1 vccd1 vccd1 _05091_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08850_ _09234_/A0 _11283_/Q _08850_/S vssd1 vssd1 vccd1 vccd1 _08851_/B sky130_fd_sc_hd__mux2_1
XFILLER_135_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07801_ _09182_/A0 _10708_/Q _09200_/S vssd1 vssd1 vccd1 vccd1 _07802_/B sky130_fd_sc_hd__mux2_1
XFILLER_112_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08781_ _08781_/A _08781_/B vssd1 vssd1 vccd1 vccd1 _11246_/D sky130_fd_sc_hd__or2_1
X_05993_ _11222_/Q _06470_/A2 _05991_/X _05992_/X vssd1 vssd1 vccd1 vccd1 _05993_/X
+ sky130_fd_sc_hd__o211a_1
X_07732_ _10667_/Q _07750_/B vssd1 vssd1 vccd1 vccd1 _07732_/X sky130_fd_sc_hd__or2_1
XFILLER_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07663_ _10626_/Q _07104_/A _07663_/S vssd1 vssd1 vccd1 vccd1 _07664_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09402_ _10214_/Q _09447_/B vssd1 vssd1 vccd1 vccd1 _11568_/D sky130_fd_sc_hd__and2_1
XFILLER_20_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06614_ _11327_/Q _10086_/A _10136_/A _11299_/Q _08243_/B vssd1 vssd1 vccd1 vccd1
+ _06614_/X sky130_fd_sc_hd__a221o_1
X_07594_ _07922_/A _07594_/B vssd1 vssd1 vccd1 vccd1 _10580_/D sky130_fd_sc_hd__or2_1
XFILLER_20_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09333_ _09985_/A1 _09343_/B _08851_/A vssd1 vssd1 vccd1 vccd1 _09333_/X sky130_fd_sc_hd__a21o_1
XFILLER_55_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06545_ _10858_/Q _06631_/A2 _06543_/X _06544_/X vssd1 vssd1 vccd1 vccd1 _06545_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09264_ _11485_/Q _09266_/B vssd1 vssd1 vccd1 vccd1 _09264_/X sky130_fd_sc_hd__or2_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06476_ _10775_/Q _06646_/A2 _08971_/A _10565_/Q vssd1 vssd1 vccd1 vccd1 _06476_/X
+ sky130_fd_sc_hd__a22o_1
X_08215_ _10942_/Q _08902_/C vssd1 vssd1 vccd1 vccd1 _08215_/X sky130_fd_sc_hd__or2_1
X_05427_ _10646_/Q _10645_/Q _05427_/S vssd1 vssd1 vccd1 vccd1 _05428_/D sky130_fd_sc_hd__mux2_1
X_09195_ _11442_/Q _09190_/Y _09193_/Y _07022_/X vssd1 vssd1 vccd1 vccd1 _11442_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08146_ _08838_/A0 _10899_/Q _08146_/S vssd1 vssd1 vccd1 vccd1 _08147_/B sky130_fd_sc_hd__mux2_1
XFILLER_140_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05358_ _11274_/Q _11273_/Q _05430_/S vssd1 vssd1 vccd1 vccd1 _05362_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08077_ _10864_/Q _08085_/B vssd1 vssd1 vccd1 vccd1 _08077_/X sky130_fd_sc_hd__or2_1
XFILLER_150_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05289_ _11172_/Q _10888_/Q _11594_/Q vssd1 vssd1 vccd1 vccd1 _05290_/D sky130_fd_sc_hd__mux2_1
XFILLER_122_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07028_ _07028_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _07241_/B sky130_fd_sc_hd__and2_1
XFILLER_134_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08979_ _09090_/A1 _08989_/B _09129_/B1 vssd1 vssd1 vccd1 vccd1 _08979_/X sky130_fd_sc_hd__a21o_1
XFILLER_76_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10941_ _11023_/CLK _10941_/D vssd1 vssd1 vccd1 vccd1 _10941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10872_ _11633_/CLK _10872_/D vssd1 vssd1 vccd1 vccd1 _10872_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11424_ _11431_/CLK _11424_/D vssd1 vssd1 vccd1 vccd1 _11424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_8 _05734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11355_ _11607_/CLK _11355_/D vssd1 vssd1 vccd1 vccd1 _11355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10306_ _11776_/CLK _10306_/D vssd1 vssd1 vccd1 vccd1 _10306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11286_ _11393_/CLK _11286_/D vssd1 vssd1 vccd1 vccd1 _11286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10237_ _11702_/CLK _10237_/D vssd1 vssd1 vccd1 vccd1 _10237_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_117_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1020 _09289_/A1 vssd1 vssd1 vccd1 vccd1 _09172_/A1 sky130_fd_sc_hd__buf_6
Xfanout1031 _08092_/A vssd1 vssd1 vccd1 vccd1 _10150_/A1 sky130_fd_sc_hd__buf_6
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1042 _10019_/A0 vssd1 vssd1 vccd1 vccd1 _09283_/A1 sky130_fd_sc_hd__buf_6
X_10168_ _10168_/A1 _10176_/B _08618_/A vssd1 vssd1 vccd1 vccd1 _10168_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1053 input112/X vssd1 vssd1 vccd1 vccd1 _10017_/A0 sky130_fd_sc_hd__buf_6
Xfanout1064 _08579_/A0 vssd1 vssd1 vccd1 vccd1 _10183_/A0 sky130_fd_sc_hd__buf_2
XFILLER_0_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1075 input102/X vssd1 vssd1 vccd1 vccd1 _10051_/A1 sky130_fd_sc_hd__buf_6
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10099_ _10149_/A1 _10087_/X _10098_/X _10155_/C1 vssd1 vssd1 vccd1 vccd1 _11751_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_63_wb_clk_i clkbuf_leaf_69_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11685_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_130_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06330_ _10846_/Q _06643_/A2 _06640_/B1 _11139_/Q _06329_/X vssd1 vssd1 vccd1 vccd1
+ _06330_/X sky130_fd_sc_hd__o221a_1
XFILLER_124_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06261_ _06257_/X _06260_/X _07083_/A _06255_/X vssd1 vssd1 vccd1 vccd1 _06261_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_129_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08000_ _08833_/A _08000_/B vssd1 vssd1 vccd1 vccd1 _10824_/D sky130_fd_sc_hd__or2_1
X_05212_ _10908_/Q _10907_/Q _05471_/A vssd1 vssd1 vccd1 vccd1 _05213_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06192_ _10400_/Q _07254_/A _07540_/A _10560_/Q vssd1 vssd1 vccd1 vccd1 _06192_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05143_ _11188_/Q _11187_/Q _05471_/A vssd1 vssd1 vccd1 vccd1 _05145_/C sky130_fd_sc_hd__mux2_1
XFILLER_116_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09951_ _10375_/Q _09567_/A _09571_/C _10694_/Q _09946_/X vssd1 vssd1 vccd1 vccd1
+ _09955_/A sky130_fd_sc_hd__a221o_1
X_05074_ _11629_/Q vssd1 vssd1 vccd1 vccd1 _05074_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08902_ _11311_/Q _08902_/B _08902_/C vssd1 vssd1 vccd1 vccd1 _08902_/X sky130_fd_sc_hd__or3_1
XFILLER_83_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09882_ _11401_/Q _09572_/A _09882_/B1 _10576_/Q vssd1 vssd1 vccd1 vccd1 _09882_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _08833_/A _08833_/B vssd1 vssd1 vccd1 vccd1 _11274_/D sky130_fd_sc_hd__or2_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08765_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08804_/B sky130_fd_sc_hd__nor2_8
XFILLER_22_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05976_ _11453_/Q _06799_/A2 _06999_/A _10341_/Q _06651_/C1 vssd1 vssd1 vccd1 vccd1
+ _05976_/X sky130_fd_sc_hd__o221a_1
Xwrapped_tms1x00_1107 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1107/HI io_oeb[37] sky130_fd_sc_hd__conb_1
XFILLER_22_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07715_ _10019_/A0 _07751_/A2 _07714_/X _07884_/C1 vssd1 vssd1 vccd1 vccd1 _10658_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1118 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1118/HI io_out[34] sky130_fd_sc_hd__conb_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1129 vssd1 vssd1 vccd1 vccd1 io_oeb[6] wrapped_tms1x00_1129/LO sky130_fd_sc_hd__conb_1
X_08695_ _08883_/A1 _11202_/Q _08695_/S vssd1 vssd1 vccd1 vccd1 _08696_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07646_ _10610_/Q _07088_/X _07651_/S vssd1 vssd1 vccd1 vccd1 _10610_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07577_ _07031_/A _10572_/Q _07593_/S vssd1 vssd1 vccd1 vccd1 _07578_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09316_ _10110_/A0 _11509_/Q _09324_/S vssd1 vssd1 vccd1 vccd1 _11509_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06528_ _11045_/Q _09059_/A _08971_/A _10967_/Q vssd1 vssd1 vccd1 vccd1 _06528_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09247_ _11477_/Q _09226_/Y _09229_/Y _07043_/X vssd1 vssd1 vccd1 vccd1 _11477_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06459_ _10944_/Q _06459_/A2 _06459_/B1 _11020_/Q vssd1 vssd1 vccd1 vccd1 _06459_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_107_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09178_ _11433_/Q _09175_/Y _09176_/Y _07227_/X vssd1 vssd1 vccd1 vccd1 _11433_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ _09395_/A0 _08140_/S _08128_/X _08841_/C1 vssd1 vssd1 vccd1 vccd1 _10890_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11140_ _11140_/CLK _11140_/D vssd1 vssd1 vccd1 vccd1 _11140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11071_ _11177_/CLK _11071_/D vssd1 vssd1 vccd1 vccd1 _11071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput101 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 input101/X sky130_fd_sc_hd__clkbuf_4
XFILLER_118_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput112 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 input112/X sky130_fd_sc_hd__buf_6
X_10022_ _10056_/A _10022_/B vssd1 vssd1 vccd1 vccd1 _11701_/D sky130_fd_sc_hd__or2_1
XFILLER_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ _11780_/CLK _10924_/D vssd1 vssd1 vccd1 vccd1 _10924_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10855_ _11269_/CLK _10855_/D vssd1 vssd1 vccd1 vccd1 _10855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _11477_/CLK _10786_/D vssd1 vssd1 vccd1 vccd1 _10786_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_110_wb_clk_i clkbuf_4_10__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10769_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ _11410_/CLK _11407_/D vssd1 vssd1 vccd1 vccd1 _11407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11338_ _11675_/CLK _11338_/D vssd1 vssd1 vccd1 vccd1 _11338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11269_ _11269_/CLK _11269_/D vssd1 vssd1 vccd1 vccd1 _11269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05830_ _11380_/Q _09060_/A _08972_/A _11340_/Q _05829_/X vssd1 vssd1 vccd1 vccd1
+ _05830_/X sky130_fd_sc_hd__o221a_1
XFILLER_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05761_ _11379_/Q _08383_/A _05757_/X _05760_/X vssd1 vssd1 vccd1 vccd1 _05762_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07500_ _10017_/A0 _07513_/S _07499_/X _07894_/C1 vssd1 vssd1 vccd1 vccd1 _10534_/D
+ sky130_fd_sc_hd__o211a_1
X_08480_ _09256_/A1 _08501_/S _08479_/X _09036_/C1 vssd1 vssd1 vccd1 vccd1 _11090_/D
+ sky130_fd_sc_hd__o211a_1
X_05692_ _05692_/A _05692_/B _05692_/C vssd1 vssd1 vccd1 vccd1 _05692_/X sky130_fd_sc_hd__or3_4
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07431_ _07141_/A _10492_/Q _07437_/S vssd1 vssd1 vccd1 vccd1 _07432_/B sky130_fd_sc_hd__mux2_1
X_07362_ _07100_/X _10453_/Q _07363_/S vssd1 vssd1 vccd1 vccd1 _10453_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09101_ _09101_/A1 _09099_/B _08873_/A vssd1 vssd1 vccd1 vccd1 _09101_/X sky130_fd_sc_hd__a21o_1
X_06313_ _11197_/Q _08668_/A _09110_/A _11247_/Q vssd1 vssd1 vccd1 vccd1 _06313_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07293_ _10415_/Q _09175_/B vssd1 vssd1 vccd1 vccd1 _07293_/X sky130_fd_sc_hd__or2_1
X_09032_ _10153_/A1 _09016_/X _09031_/X _09032_/C1 vssd1 vssd1 vccd1 vccd1 _11366_/D
+ sky130_fd_sc_hd__o211a_1
X_06244_ _10343_/Q _07152_/A _06243_/X _06651_/C1 vssd1 vssd1 vccd1 vccd1 _06244_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06175_ _11395_/Q _09082_/A _09038_/A _11375_/Q _06174_/X vssd1 vssd1 vccd1 vccd1
+ _06175_/X sky130_fd_sc_hd__o221a_1
XFILLER_89_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05126_ _10928_/Q _10927_/Q _05392_/S vssd1 vssd1 vccd1 vccd1 _05129_/B sky130_fd_sc_hd__mux2_1
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout802 _10072_/A vssd1 vssd1 vccd1 vccd1 _06632_/A2 sky130_fd_sc_hd__buf_4
X_09934_ _11664_/Q _09851_/Y _09889_/Y input8/X _09933_/Y vssd1 vssd1 vccd1 vccd1
+ _09934_/X sky130_fd_sc_hd__a221o_1
Xfanout813 _08594_/A vssd1 vssd1 vccd1 vccd1 _09977_/A sky130_fd_sc_hd__buf_4
Xfanout824 _06470_/A2 vssd1 vssd1 vccd1 vccd1 _06514_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout835 _05953_/A2 vssd1 vssd1 vccd1 vccd1 _09016_/A sky130_fd_sc_hd__buf_4
XFILLER_113_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout846 _05743_/X vssd1 vssd1 vccd1 vccd1 fanout846/X sky130_fd_sc_hd__buf_12
X_09865_ _11450_/Q _09953_/B1 _09882_/B1 _10714_/Q _09852_/X vssd1 vssd1 vccd1 vccd1
+ _09868_/C sky130_fd_sc_hd__a221o_1
Xfanout857 _06230_/A2 vssd1 vssd1 vccd1 vccd1 _06459_/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout868 _06455_/A2 vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__buf_6
Xfanout879 _07202_/A vssd1 vssd1 vccd1 vccd1 _06634_/B1 sky130_fd_sc_hd__buf_4
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08816_ _08816_/A _08816_/B vssd1 vssd1 vccd1 vccd1 _11265_/D sky130_fd_sc_hd__or2_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09796_ _11652_/Q _09771_/Y _09795_/X _09554_/B _09406_/B vssd1 vssd1 vccd1 vccd1
+ _09796_/X sky130_fd_sc_hd__o221a_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08747_ _07107_/A _08748_/S _08746_/X _08578_/A vssd1 vssd1 vccd1 vccd1 _11230_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05959_ _11382_/Q _09060_/A _09110_/A _11405_/Q _05958_/X vssd1 vssd1 vccd1 vccd1
+ _05959_/X sky130_fd_sc_hd__o221a_1
XFILLER_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _08771_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _11193_/D sky130_fd_sc_hd__or2_1
XFILLER_42_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _08649_/A _08560_/C _07847_/C vssd1 vssd1 vccd1 vccd1 _07630_/B sky130_fd_sc_hd__and3_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10640_ _10644_/CLK _10640_/D vssd1 vssd1 vccd1 vccd1 _10640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10571_ _10782_/CLK _10571_/D vssd1 vssd1 vccd1 vccd1 _10571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11123_ _11766_/CLK _11123_/D vssd1 vssd1 vccd1 vccd1 _11123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11054_ _11269_/CLK _11054_/D vssd1 vssd1 vccd1 vccd1 _11054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10005_ _10115_/A0 _11692_/Q _10008_/S vssd1 vssd1 vccd1 vccd1 _11692_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10907_ _11527_/CLK _10907_/D vssd1 vssd1 vccd1 vccd1 _10907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10838_ _11243_/CLK _10838_/D vssd1 vssd1 vccd1 vccd1 _10838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10769_ _10769_/CLK _10769_/D vssd1 vssd1 vccd1 vccd1 _10769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07980_ _10814_/Q _07015_/A _07991_/S vssd1 vssd1 vccd1 vccd1 _07981_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06931_ _10150_/A1 _10209_/Q _06934_/S vssd1 vssd1 vccd1 vccd1 _10209_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09650_ _09650_/A _09650_/B _09650_/C _09650_/D vssd1 vssd1 vccd1 vccd1 _09650_/X
+ sky130_fd_sc_hd__or4_2
X_06862_ _11462_/Q _06862_/A2 _06875_/B1 _10680_/Q vssd1 vssd1 vccd1 vccd1 _06862_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_45_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08601_ _09090_/A1 _11155_/Q _08621_/S vssd1 vssd1 vccd1 vccd1 _08602_/B sky130_fd_sc_hd__mux2_1
XFILLER_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05813_ _05805_/X _05807_/X _05812_/X _06633_/A vssd1 vssd1 vccd1 vccd1 _05813_/X
+ sky130_fd_sc_hd__a211o_1
X_09581_ _10519_/Q _09872_/A2 _09882_/B1 _10518_/Q _09577_/X vssd1 vssd1 vccd1 vccd1
+ _09586_/A sky130_fd_sc_hd__a221o_4
X_06793_ _10353_/Q _07152_/A _07455_/A _10676_/Q _06792_/X vssd1 vssd1 vccd1 vccd1
+ _06793_/X sky130_fd_sc_hd__o221a_1
XFILLER_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08532_ _08793_/A _08532_/B vssd1 vssd1 vccd1 vccd1 _11115_/D sky130_fd_sc_hd__or2_1
X_05744_ _05751_/A _05749_/A _05751_/B vssd1 vssd1 vccd1 vccd1 _05744_/Y sky130_fd_sc_hd__nor3b_4
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08463_ _11082_/Q _08467_/S _08287_/Y _07098_/B vssd1 vssd1 vccd1 vccd1 _11082_/D
+ sky130_fd_sc_hd__o22a_1
X_05675_ _11195_/Q _05537_/Y _05573_/Y _11198_/Q _05674_/X vssd1 vssd1 vccd1 vccd1
+ _05680_/B sky130_fd_sc_hd__a221o_1
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07414_ _07420_/A _07414_/B vssd1 vssd1 vccd1 vccd1 _10483_/D sky130_fd_sc_hd__or2_1
XFILLER_23_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08394_ _09283_/A1 _11038_/Q _08404_/S vssd1 vssd1 vccd1 vccd1 _08395_/B sky130_fd_sc_hd__mux2_1
XFILLER_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07345_ _10441_/Q _07350_/S _07346_/B1 _07095_/B vssd1 vssd1 vccd1 vccd1 _10441_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07276_ _07934_/A _07276_/B vssd1 vssd1 vccd1 vccd1 _10406_/D sky130_fd_sc_hd__or2_1
XFILLER_104_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09015_ _10086_/A _09015_/B _10158_/B vssd1 vssd1 vccd1 vccd1 _09035_/B sky130_fd_sc_hd__and3_4
X_06227_ _11693_/Q _06227_/A2 _10072_/A _11740_/Q _06344_/C1 vssd1 vssd1 vccd1 vccd1
+ _06227_/X sky130_fd_sc_hd__o221a_1
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06158_ _10871_/Q _06415_/A2 _06628_/B1 _10989_/Q vssd1 vssd1 vccd1 vccd1 _06158_/X
+ sky130_fd_sc_hd__o22a_1
X_05109_ _11266_/Q _11265_/Q _05397_/S vssd1 vssd1 vccd1 vccd1 _05112_/B sky130_fd_sc_hd__mux2_1
XFILLER_137_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06089_ _11493_/Q _08907_/A _08855_/A _11417_/Q vssd1 vssd1 vccd1 vccd1 _06089_/X
+ sky130_fd_sc_hd__o22a_1
Xfanout610 _06228_/A2 vssd1 vssd1 vccd1 vccd1 _09391_/A sky130_fd_sc_hd__buf_4
Xfanout621 _05737_/X vssd1 vssd1 vccd1 vccd1 _06748_/A2 sky130_fd_sc_hd__buf_8
XFILLER_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09917_ _09917_/A _09917_/B _09917_/C _09917_/D vssd1 vssd1 vccd1 vccd1 _09925_/A
+ sky130_fd_sc_hd__or4_2
Xfanout632 _09678_/A vssd1 vssd1 vccd1 vccd1 _09478_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout643 _05077_/Y vssd1 vssd1 vccd1 vccd1 _05619_/B2 sky130_fd_sc_hd__buf_8
XFILLER_28_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout654 _11655_/Q vssd1 vssd1 vccd1 vccd1 _09511_/C sky130_fd_sc_hd__clkbuf_4
Xfanout665 _05606_/B2 vssd1 vssd1 vccd1 vccd1 _05079_/A sky130_fd_sc_hd__buf_12
XFILLER_101_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout676 _11600_/Q vssd1 vssd1 vccd1 vccd1 _05349_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09848_ _10784_/Q _09882_/B1 _09567_/D _10779_/Q vssd1 vssd1 vccd1 vccd1 _09848_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout687 _05326_/S vssd1 vssd1 vccd1 vccd1 _05392_/S sky130_fd_sc_hd__buf_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout698 _06967_/A vssd1 vssd1 vccd1 vccd1 _06939_/A sky130_fd_sc_hd__buf_8
XFILLER_111_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09779_ _05429_/S _09672_/B _09674_/A _11589_/Q vssd1 vssd1 vccd1 vccd1 _09779_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11810_/CLK _11810_/D vssd1 vssd1 vccd1 vccd1 _11810_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11765_/CLK _11741_/D vssd1 vssd1 vccd1 vccd1 _11741_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11763_/CLK _11672_/D vssd1 vssd1 vccd1 vccd1 _11672_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10623_ _10798_/CLK _10623_/D vssd1 vssd1 vccd1 vccd1 _10623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ _11573_/CLK _10554_/D vssd1 vssd1 vccd1 vccd1 _10554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10485_ _10725_/CLK _10485_/D vssd1 vssd1 vccd1 vccd1 _10485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11106_ _11385_/CLK _11106_/D vssd1 vssd1 vccd1 vccd1 _11106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11037_ _11251_/CLK _11037_/D vssd1 vssd1 vccd1 vccd1 _11037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05460_ _10806_/Q _09876_/B1 _09571_/C _10764_/Q vssd1 vssd1 vccd1 vccd1 _05460_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05391_ _10743_/Q _10742_/Q _05391_/S vssd1 vssd1 vccd1 vccd1 _05395_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07130_ _10325_/Q _07145_/B vssd1 vssd1 vccd1 vccd1 _07130_/X sky130_fd_sc_hd__or2_1
XFILLER_119_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07061_ _07061_/A _10028_/A vssd1 vssd1 vccd1 vccd1 _07318_/B sky130_fd_sc_hd__and2_4
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput202 _05479_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_4
X_06012_ _06633_/A _06005_/X _06010_/X _06619_/A1 _06000_/X vssd1 vssd1 vccd1 vccd1
+ _06012_/X sky130_fd_sc_hd__o311a_1
XFILLER_86_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07963_ _07052_/X _07883_/B _07962_/X vssd1 vssd1 vccd1 vccd1 _10804_/D sky130_fd_sc_hd__a21o_1
XFILLER_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06914_ _10149_/A1 _06922_/B _08664_/A vssd1 vssd1 vccd1 vccd1 _06914_/X sky130_fd_sc_hd__a21o_1
X_09702_ _11638_/Q _11642_/Q _09702_/S vssd1 vssd1 vccd1 vccd1 _09703_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07894_ _07076_/A _07970_/S _07893_/X _07894_/C1 vssd1 vssd1 vccd1 vccd1 _10765_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06845_ _11461_/Q _06875_/A2 _06844_/X _06878_/C1 vssd1 vssd1 vccd1 vccd1 _06845_/X
+ sky130_fd_sc_hd__o211a_1
X_09633_ _09633_/A _09633_/B _09633_/C _09633_/D vssd1 vssd1 vccd1 vccd1 _09636_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09564_ _09564_/A _09564_/B vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__nor2_4
X_06776_ _10412_/Q _07254_/A vssd1 vssd1 vccd1 vccd1 _06776_/X sky130_fd_sc_hd__or2_1
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08515_ _11107_/Q _08545_/B vssd1 vssd1 vccd1 vccd1 _08515_/X sky130_fd_sc_hd__or2_1
X_05727_ _05727_/A _05727_/B _05727_/C _05727_/D vssd1 vssd1 vccd1 vccd1 _05728_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_110_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09495_ _09528_/A _09500_/B _09495_/C vssd1 vssd1 vccd1 vccd1 _09496_/A sky130_fd_sc_hd__nand3_1
XFILLER_145_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08446_ _11067_/Q _08436_/Y _08439_/Y _07333_/X vssd1 vssd1 vccd1 vccd1 _11067_/D
+ sky130_fd_sc_hd__a22o_1
X_05658_ _11247_/Q _05549_/Y _05603_/Y _11243_/Q vssd1 vssd1 vccd1 vccd1 _05661_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08377_ _08757_/A _08377_/B vssd1 vssd1 vccd1 vccd1 _11030_/D sky130_fd_sc_hd__or2_1
X_05589_ _05631_/A2 _10202_/Q _10198_/Q _05631_/B1 _05587_/X vssd1 vssd1 vccd1 vccd1
+ _05589_/X sky130_fd_sc_hd__a221o_1
XFILLER_17_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07328_ _10428_/Q _07322_/Y _07326_/Y _07008_/X vssd1 vssd1 vccd1 vccd1 _10428_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07259_ _10017_/A0 _10398_/Q _07259_/S vssd1 vssd1 vccd1 vccd1 _07260_/B sky130_fd_sc_hd__mux2_1
XFILLER_104_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10270_ _11703_/CLK _10270_/D vssd1 vssd1 vccd1 vccd1 _10270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout440 _05204_/X vssd1 vssd1 vccd1 vccd1 _09566_/A sky130_fd_sc_hd__buf_8
XFILLER_63_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout451 _05146_/Y vssd1 vssd1 vccd1 vccd1 _09877_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout462 _07018_/B vssd1 vssd1 vccd1 vccd1 _07107_/B sky130_fd_sc_hd__buf_8
Xfanout473 _06996_/C1 vssd1 vssd1 vccd1 vccd1 _06990_/C1 sky130_fd_sc_hd__buf_4
XFILLER_24_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout484 _07882_/C1 vssd1 vssd1 vccd1 vccd1 _09201_/A1 sky130_fd_sc_hd__buf_6
XFILLER_74_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout495 _09993_/C1 vssd1 vssd1 vccd1 vccd1 _10177_/C1 sky130_fd_sc_hd__buf_2
XFILLER_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _11735_/CLK _11724_/D vssd1 vssd1 vccd1 vccd1 _11724_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11655_ _11663_/CLK _11655_/D vssd1 vssd1 vccd1 vccd1 _11655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ _11262_/CLK _10606_/D vssd1 vssd1 vccd1 vccd1 _10606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_88_wb_clk_i clkbuf_leaf_88_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11657_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11586_ _11652_/CLK _11586_/D vssd1 vssd1 vccd1 vccd1 _11586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10537_ _11442_/CLK _10537_/D vssd1 vssd1 vccd1 vccd1 _10537_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11307_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10468_ _11140_/CLK _10468_/D vssd1 vssd1 vccd1 vccd1 _10468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10399_ _10785_/CLK _10399_/D vssd1 vssd1 vccd1 vccd1 _10399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06630_ _10948_/Q _06630_/A2 _06630_/B1 _11024_/Q vssd1 vssd1 vccd1 vccd1 _06630_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06561_ _10405_/Q _06645_/A2 _09109_/A _10542_/Q vssd1 vssd1 vccd1 vccd1 _06561_/X
+ sky130_fd_sc_hd__a22o_1
X_08300_ _08300_/A _08665_/C _09038_/C vssd1 vssd1 vccd1 vccd1 _08832_/S sky130_fd_sc_hd__or3_4
X_05512_ input5/X _11338_/Q _10213_/Q vssd1 vssd1 vccd1 vccd1 _11608_/D sky130_fd_sc_hd__mux2_1
X_09280_ _09280_/A1 _09288_/B _09290_/B1 vssd1 vssd1 vccd1 vccd1 _09280_/X sky130_fd_sc_hd__a21o_1
X_06492_ _06663_/A _10233_/Q vssd1 vssd1 vccd1 vccd1 _06493_/B sky130_fd_sc_hd__and2_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08231_ _10949_/Q _08324_/B vssd1 vssd1 vccd1 vccd1 _08231_/X sky130_fd_sc_hd__or2_1
X_05443_ _10681_/Q _09953_/B1 _09565_/B _10665_/Q _05442_/X vssd1 vssd1 vccd1 vccd1
+ _05451_/C sky130_fd_sc_hd__a221o_1
XFILLER_53_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08162_ _08760_/A0 _10907_/Q _08162_/S vssd1 vssd1 vccd1 vccd1 _08163_/B sky130_fd_sc_hd__mux2_1
X_05374_ _10870_/Q _10869_/Q _05427_/S vssd1 vssd1 vccd1 vccd1 _05378_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07113_ _10310_/Q _07126_/B _07186_/S _07324_/B vssd1 vssd1 vccd1 vccd1 _10310_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_88_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08093_ _08015_/S _08092_/X _08091_/X _08427_/A vssd1 vssd1 vccd1 vccd1 _10871_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_1348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07044_ _10279_/Q _07043_/X _07044_/S vssd1 vssd1 vccd1 vccd1 _10279_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08995_ _11349_/Q _09013_/B vssd1 vssd1 vccd1 vccd1 _08995_/X sky130_fd_sc_hd__or2_1
XFILLER_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07946_ _10788_/Q _07941_/Y _07944_/Y _07227_/X vssd1 vssd1 vccd1 vccd1 _10788_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07877_ _10757_/Q _07893_/B vssd1 vssd1 vccd1 vccd1 _07877_/X sky130_fd_sc_hd__or2_1
X_09616_ _10387_/Q _09944_/B1 _09947_/B1 _10391_/Q _09603_/X vssd1 vssd1 vccd1 vccd1
+ _09617_/D sky130_fd_sc_hd__a221o_1
X_06828_ _10334_/Q _06856_/A2 _06685_/B _11721_/Q vssd1 vssd1 vccd1 vccd1 _06828_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06759_ _10296_/Q _07046_/A _07190_/A _10491_/Q _06758_/X vssd1 vssd1 vccd1 vccd1
+ _06759_/X sky130_fd_sc_hd__o221a_1
X_09547_ _11664_/Q _09538_/X _09542_/X vssd1 vssd1 vccd1 vccd1 _09547_/X sky130_fd_sc_hd__a21o_1
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09478_ _09478_/A _09554_/A _09478_/C vssd1 vssd1 vccd1 vccd1 _11602_/D sky130_fd_sc_hd__and3_1
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08429_ _11054_/Q _08425_/Y _08426_/Y _08441_/B2 vssd1 vssd1 vccd1 vccd1 _11054_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_156_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11440_ _11473_/CLK _11440_/D vssd1 vssd1 vccd1 vccd1 _11440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11371_ _11431_/CLK _11371_/D vssd1 vssd1 vccd1 vccd1 _11371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10322_ _10727_/CLK _10322_/D vssd1 vssd1 vccd1 vccd1 _10322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10253_ _11712_/CLK _10253_/D vssd1 vssd1 vccd1 vccd1 _10253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10184_ _10184_/A0 _11805_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _11805_/D sky130_fd_sc_hd__mux2_1
XFILLER_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_135_wb_clk_i clkbuf_4_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11716_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout270 _08200_/X vssd1 vssd1 vccd1 vccd1 _08225_/S sky130_fd_sc_hd__clkbuf_8
Xfanout281 _09206_/B vssd1 vssd1 vccd1 vccd1 _09218_/S sky130_fd_sc_hd__buf_8
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout292 _07819_/Y vssd1 vssd1 vccd1 vccd1 _07839_/A2 sky130_fd_sc_hd__buf_8
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11707_ _11716_/CLK _11707_/D vssd1 vssd1 vccd1 vccd1 _11707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11638_ _11652_/CLK _11638_/D vssd1 vssd1 vccd1 vccd1 _11638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11569_ _11573_/CLK _11569_/D vssd1 vssd1 vccd1 vccd1 _11569_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05090_ _10954_/Q vssd1 vssd1 vccd1 vccd1 _08241_/A sky130_fd_sc_hd__inv_2
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07800_ _07818_/A _07800_/B vssd1 vssd1 vccd1 vccd1 _10707_/D sky130_fd_sc_hd__or2_1
X_08780_ _08987_/A1 _11246_/Q _08802_/S vssd1 vssd1 vccd1 vccd1 _08781_/B sky130_fd_sc_hd__mux2_1
X_05992_ _10463_/Q _06642_/A2 _08469_/B _10978_/Q vssd1 vssd1 vccd1 vccd1 _05992_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07731_ _08883_/A1 _07751_/A2 _07730_/X _07894_/C1 vssd1 vssd1 vccd1 vccd1 _10666_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07662_ _10625_/Q _07663_/S _07233_/S _07318_/B vssd1 vssd1 vccd1 vccd1 _10625_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09401_ _10190_/A0 _11567_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _11567_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06613_ _11047_/Q _05736_/Y _05746_/X _10969_/Q vssd1 vssd1 vccd1 vccd1 _06613_/X
+ sky130_fd_sc_hd__a22o_1
X_07593_ _07036_/A _10580_/Q _07593_/S vssd1 vssd1 vccd1 vccd1 _07594_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06544_ _10946_/Q _06630_/A2 _06630_/B1 _11022_/Q vssd1 vssd1 vccd1 vccd1 _06544_/X
+ sky130_fd_sc_hd__o22a_1
X_09332_ _09364_/A1 _09326_/X _09331_/X _09993_/C1 vssd1 vssd1 vccd1 vccd1 _11520_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09263_ _11484_/Q _09249_/X _09262_/X vssd1 vssd1 vccd1 vccd1 _11484_/D sky130_fd_sc_hd__a21o_1
XFILLER_21_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06475_ _10404_/Q _06645_/A2 _09131_/A _10664_/Q vssd1 vssd1 vccd1 vccd1 _06475_/X
+ sky130_fd_sc_hd__a22o_1
X_08214_ _08839_/A _08214_/B vssd1 vssd1 vccd1 vccd1 _10941_/D sky130_fd_sc_hd__or2_1
X_05426_ _10649_/Q _10648_/Q _05426_/S vssd1 vssd1 vccd1 vccd1 _05428_/C sky130_fd_sc_hd__mux2_1
XFILLER_18_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09194_ _11441_/Q _09190_/Y _09193_/Y _07019_/X vssd1 vssd1 vccd1 vccd1 _11441_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08145_ _07107_/A _08140_/S _08144_/X _08841_/C1 vssd1 vssd1 vccd1 vccd1 _10898_/D
+ sky130_fd_sc_hd__o211a_1
X_05357_ _05357_/A _05357_/B vssd1 vssd1 vccd1 vccd1 _05357_/Y sky130_fd_sc_hd__nor2_8
XFILLER_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08076_ _09141_/A1 _08083_/S _08075_/X _08753_/C1 vssd1 vssd1 vccd1 vccd1 _10863_/D
+ sky130_fd_sc_hd__o211a_1
X_05288_ _10892_/Q _10891_/Q _05372_/S vssd1 vssd1 vccd1 vccd1 _05290_/C sky130_fd_sc_hd__mux2_1
XFILLER_134_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07027_ _10273_/Q _07026_/X _07038_/S vssd1 vssd1 vccd1 vccd1 _10273_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08978_ _09276_/A1 _08972_/X _08977_/X _09122_/C1 vssd1 vssd1 vccd1 vccd1 _11341_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07929_ _08423_/A1 _10782_/Q _09218_/S vssd1 vssd1 vccd1 vccd1 _07930_/B sky130_fd_sc_hd__mux2_1
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10940_ _11312_/CLK _10940_/D vssd1 vssd1 vccd1 vccd1 _10940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10871_ _11634_/CLK _10871_/D vssd1 vssd1 vccd1 vccd1 _10871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11423_ _11431_/CLK _11423_/D vssd1 vssd1 vccd1 vccd1 _11423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_9 _05734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ _11607_/CLK _11354_/D vssd1 vssd1 vccd1 vccd1 _11354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10305_ _11780_/CLK _10305_/D vssd1 vssd1 vccd1 vccd1 _10305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11285_ _11411_/CLK _11285_/D vssd1 vssd1 vccd1 vccd1 _11285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10236_ _11233_/CLK _10236_/D vssd1 vssd1 vccd1 vccd1 _10236_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1010 input117/X vssd1 vssd1 vccd1 vccd1 _07057_/A sky130_fd_sc_hd__buf_12
XFILLER_105_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1021 _10177_/A1 vssd1 vssd1 vccd1 vccd1 _09289_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_67_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10167_ _11795_/Q _10159_/X _10166_/X vssd1 vssd1 vccd1 vccd1 _11795_/D sky130_fd_sc_hd__a21o_1
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1032 input114/X vssd1 vssd1 vccd1 vccd1 _08092_/A sky130_fd_sc_hd__buf_6
Xfanout1043 _10019_/A0 vssd1 vssd1 vccd1 vccd1 _10171_/A1 sky130_fd_sc_hd__buf_6
XFILLER_48_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1054 _09395_/A0 vssd1 vssd1 vccd1 vccd1 _10112_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1065 _10142_/A1 vssd1 vssd1 vccd1 vccd1 _08579_/A0 sky130_fd_sc_hd__buf_4
Xfanout1076 input102/X vssd1 vssd1 vccd1 vccd1 _07933_/A0 sky130_fd_sc_hd__clkbuf_2
X_10098_ _11751_/Q _10104_/B vssd1 vssd1 vccd1 vccd1 _10098_/X sky130_fd_sc_hd__or2_1
XFILLER_43_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_32_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11312_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06260_ _11130_/Q _06635_/A2 _06259_/X _11869_/A vssd1 vssd1 vccd1 vccd1 _06260_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05211_ _10903_/Q _10429_/Q _08956_/B vssd1 vssd1 vccd1 vccd1 _05213_/C sky130_fd_sc_hd__mux2_1
XFILLER_128_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06191_ _10659_/Q _06806_/B1 _06728_/B1 _10536_/Q vssd1 vssd1 vccd1 vccd1 _06191_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05142_ _11186_/Q _11185_/Q _05419_/S vssd1 vssd1 vccd1 vccd1 _05145_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09950_ _10370_/Q _09565_/A _09950_/B1 _10366_/Q vssd1 vssd1 vccd1 vccd1 _09950_/X
+ sky130_fd_sc_hd__a22o_1
X_05073_ _11651_/Q vssd1 vssd1 vccd1 vccd1 _09775_/B sky130_fd_sc_hd__inv_2
XFILLER_100_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08901_ _11310_/Q _08901_/A1 _08901_/S vssd1 vssd1 vccd1 vccd1 _11310_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _10570_/Q _09881_/A2 _09881_/B1 _10560_/Q vssd1 vssd1 vccd1 vccd1 _09887_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08832_ _08970_/A1 _11274_/Q _08832_/S vssd1 vssd1 vccd1 vccd1 _08833_/B sky130_fd_sc_hd__mux2_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05975_ _10749_/Q _07853_/A vssd1 vssd1 vccd1 vccd1 _05975_/X sky130_fd_sc_hd__or2_1
X_08763_ _08665_/A _08760_/S _08762_/X _09267_/C1 vssd1 vssd1 vccd1 vccd1 _11238_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapped_tms1x00_1108 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1108/HI io_out[0] sky130_fd_sc_hd__conb_1
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07714_ _10658_/Q _07750_/B vssd1 vssd1 vccd1 vccd1 _07714_/X sky130_fd_sc_hd__or2_1
Xwrapped_tms1x00_1119 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1119/HI io_out[35] sky130_fd_sc_hd__conb_1
XFILLER_22_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _08933_/A1 _08695_/S _08693_/X _08791_/C1 vssd1 vssd1 vccd1 vccd1 _11201_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07645_ _08050_/A _07645_/B vssd1 vssd1 vccd1 vccd1 _07651_/S sky130_fd_sc_hd__or2_4
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07576_ _07930_/A _07576_/B vssd1 vssd1 vccd1 vccd1 _10571_/D sky130_fd_sc_hd__or2_1
XFILLER_0_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09315_ _09999_/A0 _11508_/Q _09324_/S vssd1 vssd1 vccd1 vccd1 _11508_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06527_ _06521_/X _06526_/X _11872_/A vssd1 vssd1 vccd1 vccd1 _06527_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _11476_/Q _09226_/Y _09229_/Y _07040_/X vssd1 vssd1 vccd1 vccd1 _11476_/D
+ sky130_fd_sc_hd__a22o_1
X_06458_ _10653_/Q _06629_/A2 _06589_/A2 _11098_/Q _07690_/B vssd1 vssd1 vccd1 vccd1
+ _06458_/X sky130_fd_sc_hd__o221a_1
XFILLER_107_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05409_ _11284_/Q _11283_/Q _06942_/A vssd1 vssd1 vccd1 vccd1 _05411_/C sky130_fd_sc_hd__mux2_1
X_09177_ _11432_/Q _09175_/Y _09176_/Y _07008_/X vssd1 vssd1 vccd1 vccd1 _11432_/D
+ sky130_fd_sc_hd__a22o_1
X_06389_ _10942_/Q _06630_/A2 _06629_/B1 _11096_/Q vssd1 vssd1 vccd1 vccd1 _06389_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08128_ _10890_/Q _08637_/C vssd1 vssd1 vccd1 vccd1 _08128_/X sky130_fd_sc_hd__or2_1
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08059_ _10855_/Q _08426_/B vssd1 vssd1 vccd1 vccd1 _08059_/X sky130_fd_sc_hd__or2_1
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11070_ _11177_/CLK _11070_/D vssd1 vssd1 vccd1 vccd1 _11070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput102 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 input102/X sky130_fd_sc_hd__clkbuf_2
X_10021_ _10021_/A0 _11701_/Q _10028_/B vssd1 vssd1 vccd1 vccd1 _10022_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput113 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 input113/X sky130_fd_sc_hd__buf_2
XFILLER_118_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10923_ _11781_/CLK _10923_/D vssd1 vssd1 vccd1 vccd1 _10923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10854_ _11604_/CLK _10854_/D vssd1 vssd1 vccd1 vccd1 _10854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _10785_/CLK _10785_/D vssd1 vssd1 vccd1 vccd1 _10785_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_125_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11406_ _11495_/CLK _11406_/D vssd1 vssd1 vccd1 vccd1 _11406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11337_ _11675_/CLK _11337_/D vssd1 vssd1 vccd1 vccd1 _11337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11268_ _11268_/CLK _11268_/D vssd1 vssd1 vccd1 vccd1 _11268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10219_ _10765_/CLK _10219_/D vssd1 vssd1 vccd1 vccd1 _10219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11199_ _11319_/CLK _11199_/D vssd1 vssd1 vccd1 vccd1 _11199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05760_ _11422_/Q _09154_/A _05759_/X _06670_/D1 vssd1 vssd1 vccd1 vccd1 _05760_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05691_ _05691_/A _05691_/B _05691_/C vssd1 vssd1 vccd1 vccd1 _05692_/C sky130_fd_sc_hd__or3_1
XFILLER_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07430_ _10050_/A _07430_/B vssd1 vssd1 vccd1 vccd1 _10491_/D sky130_fd_sc_hd__or2_1
XFILLER_39_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07361_ _08441_/B2 _10452_/Q _07363_/S vssd1 vssd1 vccd1 vccd1 _10452_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09100_ _09289_/A1 _09082_/X _09099_/X _09289_/C1 vssd1 vssd1 vccd1 vccd1 _11397_/D
+ sky130_fd_sc_hd__o211a_1
X_06312_ _11321_/Q _08907_/A _08855_/A _11293_/Q _06718_/C1 vssd1 vssd1 vccd1 vccd1
+ _06312_/X sky130_fd_sc_hd__o221a_1
X_07292_ _07812_/A _07292_/B vssd1 vssd1 vccd1 vccd1 _10414_/D sky130_fd_sc_hd__or2_1
XFILLER_31_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09031_ _11366_/Q _09035_/B vssd1 vssd1 vccd1 vccd1 _09031_/X sky130_fd_sc_hd__or2_1
X_06243_ _11441_/Q _07778_/A _06805_/B1 _10537_/Q _06242_/X vssd1 vssd1 vccd1 vccd1
+ _06243_/X sky130_fd_sc_hd__o221a_1
XFILLER_117_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06174_ _11494_/Q _08907_/A _08855_/A _11418_/Q vssd1 vssd1 vccd1 vccd1 _06174_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_89_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05125_ _10615_/Q _10614_/Q _05398_/S vssd1 vssd1 vccd1 vccd1 _05129_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09933_ _11664_/Q _09938_/B vssd1 vssd1 vccd1 vccd1 _09933_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout803 _10072_/A vssd1 vssd1 vccd1 vccd1 _06924_/A sky130_fd_sc_hd__buf_6
XFILLER_89_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout814 _06412_/B1 vssd1 vssd1 vccd1 vccd1 _08594_/A sky130_fd_sc_hd__clkbuf_8
Xfanout825 _06470_/A2 vssd1 vssd1 vccd1 vccd1 _08650_/A sky130_fd_sc_hd__buf_6
XFILLER_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout836 fanout846/X vssd1 vssd1 vccd1 vccd1 _05953_/A2 sky130_fd_sc_hd__buf_4
Xfanout847 _10086_/A vssd1 vssd1 vccd1 vccd1 _08649_/A sky130_fd_sc_hd__buf_12
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _11443_/Q _09884_/A2 _09567_/D _10709_/Q _09863_/X vssd1 vssd1 vccd1 vccd1
+ _09868_/B sky130_fd_sc_hd__a221o_1
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout858 _06540_/A2 vssd1 vssd1 vccd1 vccd1 _06976_/A sky130_fd_sc_hd__buf_6
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout869 _06455_/A2 vssd1 vssd1 vccd1 vccd1 _09154_/A sky130_fd_sc_hd__buf_4
X_08815_ _11265_/Q _10132_/A0 _08820_/S vssd1 vssd1 vccd1 vccd1 _08816_/B sky130_fd_sc_hd__mux2_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _05430_/S _09672_/B _09674_/A _11593_/Q vssd1 vssd1 vccd1 vccd1 _09795_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_100_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08746_ _11230_/Q _08750_/B vssd1 vssd1 vccd1 vccd1 _08746_/X sky130_fd_sc_hd__or2_1
X_05958_ _11491_/Q _08907_/A _08855_/A _11415_/Q vssd1 vssd1 vccd1 vccd1 _05958_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_207 _10086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05889_ _11794_/Q _10159_/A _09293_/A _11500_/Q vssd1 vssd1 vccd1 vccd1 _05889_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _09141_/A1 _11193_/Q _08695_/S vssd1 vssd1 vccd1 vccd1 _08678_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07628_ _07235_/X _10600_/Q _07628_/S vssd1 vssd1 vccd1 vccd1 _10600_/D sky130_fd_sc_hd__mux2_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07559_ _09129_/A1 _10563_/Q _07589_/S vssd1 vssd1 vccd1 vccd1 _07560_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ _10773_/CLK _10570_/D vssd1 vssd1 vccd1 vccd1 _10570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09229_ _09229_/A _09243_/C vssd1 vssd1 vccd1 vccd1 _09229_/Y sky130_fd_sc_hd__nand2_4
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11122_ _11572_/CLK _11122_/D vssd1 vssd1 vccd1 vccd1 _11122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11053_ _11269_/CLK _11053_/D vssd1 vssd1 vccd1 vccd1 _11053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10004_ _10114_/A0 _11691_/Q _10008_/S vssd1 vssd1 vccd1 vccd1 _11691_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ _11284_/CLK _10906_/D vssd1 vssd1 vccd1 vccd1 _10906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10837_ _11657_/CLK _10837_/D vssd1 vssd1 vccd1 vccd1 _10837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10768_ _11439_/CLK _10768_/D vssd1 vssd1 vccd1 vccd1 _10768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10699_ _11622_/CLK _10699_/D vssd1 vssd1 vccd1 vccd1 _10699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06930_ _10149_/A1 _10208_/Q _06934_/S vssd1 vssd1 vccd1 vccd1 _10208_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06861_ _10768_/Q _06861_/B vssd1 vssd1 vccd1 vccd1 _06861_/X sky130_fd_sc_hd__or2_1
XFILLER_95_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08600_ _08618_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _11154_/D sky130_fd_sc_hd__or2_1
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05812_ _11087_/Q _06629_/B1 _05808_/X _05811_/X vssd1 vssd1 vccd1 vccd1 _05812_/X
+ sky130_fd_sc_hd__o211a_1
X_09580_ _10267_/Q _09566_/B _09566_/C _10268_/Q vssd1 vssd1 vccd1 vccd1 _09580_/X
+ sky130_fd_sc_hd__a22o_1
X_06792_ _10808_/Q _07853_/A _07540_/A _10577_/Q vssd1 vssd1 vccd1 vccd1 _06792_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_83_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05743_ _05745_/A _05749_/A _05751_/B vssd1 vssd1 vccd1 vccd1 _05743_/X sky130_fd_sc_hd__or3_4
XFILLER_36_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08531_ _08846_/A0 _11115_/Q _08537_/S vssd1 vssd1 vccd1 vccd1 _08532_/B sky130_fd_sc_hd__mux2_1
XFILLER_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08462_ _08749_/A _08462_/B vssd1 vssd1 vccd1 vccd1 _11081_/D sky130_fd_sc_hd__or2_1
X_05674_ _11208_/Q _05518_/Y _05524_/Y _11199_/Q vssd1 vssd1 vccd1 vccd1 _05674_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07413_ _07057_/A _10483_/Q _07429_/S vssd1 vssd1 vccd1 vccd1 _07414_/B sky130_fd_sc_hd__mux2_1
X_08393_ _08771_/A _08393_/B vssd1 vssd1 vccd1 vccd1 _11037_/D sky130_fd_sc_hd__or2_1
XFILLER_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07344_ _10440_/Q _07337_/X _07346_/B1 _07617_/B vssd1 vssd1 vccd1 vccd1 _10440_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07275_ _07211_/A _10406_/Q _09187_/S vssd1 vssd1 vccd1 vccd1 _07276_/B sky130_fd_sc_hd__mux2_1
XFILLER_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06226_ _11673_/Q _09965_/A _09314_/A _11515_/Q _06225_/X vssd1 vssd1 vccd1 vccd1
+ _06226_/X sky130_fd_sc_hd__o221a_1
X_09014_ _10106_/A1 _08994_/X _09013_/X _09036_/C1 vssd1 vssd1 vccd1 vccd1 _11358_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06157_ _06153_/X _06156_/X _07083_/A _06151_/X vssd1 vssd1 vccd1 vccd1 _06157_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05108_ _10604_/Q _10603_/Q _05429_/S vssd1 vssd1 vccd1 vccd1 _05112_/A sky130_fd_sc_hd__mux2_1
X_06088_ _11394_/Q _09082_/A _08972_/A _11344_/Q vssd1 vssd1 vccd1 vccd1 _06088_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout600 _05774_/Y vssd1 vssd1 vccd1 vccd1 _07151_/B sky130_fd_sc_hd__buf_8
Xfanout611 _06228_/A2 vssd1 vssd1 vccd1 vccd1 _09965_/A sky130_fd_sc_hd__buf_6
XFILLER_63_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout622 _06696_/A2 vssd1 vssd1 vccd1 vccd1 _09326_/A sky130_fd_sc_hd__buf_4
X_09916_ _10474_/Q _09566_/A _09572_/B _10492_/Q _09915_/X vssd1 vssd1 vccd1 vccd1
+ _09917_/D sky130_fd_sc_hd__a221o_1
Xfanout633 _09447_/B vssd1 vssd1 vccd1 vccd1 _09678_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_154_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout644 _05076_/Y vssd1 vssd1 vccd1 vccd1 _05628_/A2 sky130_fd_sc_hd__buf_6
XFILLER_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout655 _11654_/Q vssd1 vssd1 vccd1 vccd1 _09515_/B sky130_fd_sc_hd__clkbuf_4
Xfanout666 _11624_/Q vssd1 vssd1 vccd1 vccd1 _05606_/B2 sky130_fd_sc_hd__buf_12
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ _10783_/Q _09879_/B1 _09877_/B1 _11456_/Q _09846_/X vssd1 vssd1 vccd1 vccd1
+ _09850_/C sky130_fd_sc_hd__a221o_1
Xfanout677 _05398_/S vssd1 vssd1 vccd1 vccd1 _05385_/S sky130_fd_sc_hd__buf_6
XFILLER_59_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout688 _05414_/S vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__buf_6
XFILLER_101_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout699 _11595_/Q vssd1 vssd1 vccd1 vccd1 _06967_/A sky130_fd_sc_hd__buf_6
XFILLER_85_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _11647_/Q _08950_/B _09773_/X _09777_/X _09407_/A vssd1 vssd1 vccd1 vccd1
+ _11647_/D sky130_fd_sc_hd__o221a_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _08745_/A _08729_/B vssd1 vssd1 vccd1 vccd1 _11221_/D sky130_fd_sc_hd__or2_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11756_/CLK _11740_/D vssd1 vssd1 vccd1 vccd1 _11740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11671_ _11763_/CLK _11671_/D vssd1 vssd1 vccd1 vccd1 _11671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10622_ _11702_/CLK _10622_/D vssd1 vssd1 vccd1 vccd1 _10622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553_ _11472_/CLK _10553_/D vssd1 vssd1 vccd1 vccd1 _10553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _11743_/CLK _10484_/D vssd1 vssd1 vccd1 vccd1 _10484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ _11428_/CLK _11105_/D vssd1 vssd1 vccd1 vccd1 _11105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11036_ _11243_/CLK _11036_/D vssd1 vssd1 vccd1 vccd1 _11036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11869_ _11869_/A vssd1 vssd1 vccd1 vccd1 _11869_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05390_ _05390_/A _05390_/B vssd1 vssd1 vccd1 vccd1 _05390_/Y sky130_fd_sc_hd__nor2_8
XFILLER_119_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07060_ _10288_/Q _07047_/B _07490_/S _07316_/B vssd1 vssd1 vccd1 vccd1 _10288_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06011_ _07151_/B _05984_/X _05989_/X _05973_/X vssd1 vssd1 vccd1 vccd1 _06011_/X
+ sky130_fd_sc_hd__a211o_2
Xoutput203 _05507_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_4
XFILLER_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07962_ _10804_/Q _09227_/A _07871_/S _09192_/A vssd1 vssd1 vccd1 vccd1 _07962_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09701_ _09703_/A _09701_/B vssd1 vssd1 vccd1 vccd1 _11641_/D sky130_fd_sc_hd__or2_1
X_06913_ _10185_/A0 _06903_/X _06912_/X _06990_/C1 vssd1 vssd1 vccd1 vccd1 _10197_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07893_ _10765_/Q _07893_/B vssd1 vssd1 vccd1 vccd1 _07893_/X sky130_fd_sc_hd__or2_1
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ _10717_/Q _09566_/A _09565_/B _10725_/Q _09628_/X vssd1 vssd1 vccd1 vccd1
+ _09633_/D sky130_fd_sc_hd__a221o_1
X_06844_ _11475_/Q _07153_/A _06877_/B1 _11399_/Q _06843_/X vssd1 vssd1 vccd1 vccd1
+ _06844_/X sky130_fd_sc_hd__o221a_1
XFILLER_56_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09563_ _11659_/Q _11644_/Q vssd1 vssd1 vccd1 vccd1 _09564_/B sky130_fd_sc_hd__nor2_1
XFILLER_110_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06775_ _10331_/Q _07539_/A _06771_/X _06774_/X vssd1 vssd1 vccd1 vccd1 _06775_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08514_ _09090_/A1 _08537_/S _08513_/X _09168_/C1 vssd1 vssd1 vccd1 vccd1 _11106_/D
+ sky130_fd_sc_hd__o211a_1
X_05726_ _10957_/Q _05531_/Y _05555_/Y _10966_/Q vssd1 vssd1 vccd1 vccd1 _05727_/D
+ sky130_fd_sc_hd__a22o_1
X_09494_ _09511_/C _09515_/C _09515_/B vssd1 vssd1 vccd1 vccd1 _09495_/C sky130_fd_sc_hd__nor3b_2
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08445_ _11066_/Q _08437_/Y _08438_/Y _07318_/X vssd1 vssd1 vccd1 vccd1 _11066_/D
+ sky130_fd_sc_hd__o22a_1
X_05657_ _11256_/Q _05543_/Y _05615_/Y _11252_/Q vssd1 vssd1 vccd1 vccd1 _05661_/A
+ sky130_fd_sc_hd__a22o_1
X_05588_ _05630_/A2 _10196_/Q _10193_/Q _05079_/A _05586_/X vssd1 vssd1 vccd1 vccd1
+ _05591_/A sky130_fd_sc_hd__a221o_4
X_08376_ _10153_/A1 _11030_/Q _08439_/B vssd1 vssd1 vccd1 vccd1 _08377_/B sky130_fd_sc_hd__mux2_1
XFILLER_149_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07327_ _10427_/Q _07322_/Y _07324_/X _07326_/Y vssd1 vssd1 vccd1 vccd1 _10427_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07258_ _07916_/A _07258_/B vssd1 vssd1 vccd1 vccd1 _10397_/D sky130_fd_sc_hd__or2_1
XFILLER_104_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06209_ _06663_/A _10228_/Q _06535_/A vssd1 vssd1 vccd1 vccd1 _06209_/X sky130_fd_sc_hd__a21o_1
X_07189_ _07190_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _07191_/B sky130_fd_sc_hd__nor2_8
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout430 _05259_/Y vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__buf_6
XFILLER_28_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout441 _05204_/X vssd1 vssd1 vccd1 vccd1 _09874_/A2 sky130_fd_sc_hd__buf_4
XFILLER_120_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout452 _05135_/Y vssd1 vssd1 vccd1 vccd1 _09570_/A sky130_fd_sc_hd__buf_8
Xfanout463 _08345_/C1 vssd1 vssd1 vccd1 vccd1 _08841_/C1 sky130_fd_sc_hd__buf_4
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout474 _10153_/C1 vssd1 vssd1 vccd1 vccd1 _06996_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout485 _07866_/C1 vssd1 vssd1 vccd1 vccd1 _07868_/C1 sky130_fd_sc_hd__buf_6
XFILLER_87_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout496 fanout510/X vssd1 vssd1 vccd1 vccd1 _09993_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_58_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11756_/CLK _11723_/D vssd1 vssd1 vccd1 vccd1 _11723_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11663_/CLK _11654_/D vssd1 vssd1 vccd1 vccd1 _11654_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ _11262_/CLK _10605_/D vssd1 vssd1 vccd1 vccd1 _10605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11585_ _11652_/CLK _11585_/D vssd1 vssd1 vccd1 vccd1 _11585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10536_ _10808_/CLK _10536_/D vssd1 vssd1 vccd1 vccd1 _10536_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_109_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10467_ _11307_/CLK _10467_/D vssd1 vssd1 vccd1 vccd1 _10467_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_57_wb_clk_i clkbuf_leaf_88_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11280_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10398_ _10805_/CLK _10398_/D vssd1 vssd1 vccd1 vccd1 _10398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11019_ _11312_/CLK _11019_/D vssd1 vssd1 vccd1 vccd1 _11019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06560_ _10777_/Q _06646_/A2 _06649_/A2 _10347_/Q _06873_/D1 vssd1 vssd1 vccd1 vccd1
+ _06560_/X sky130_fd_sc_hd__a221o_1
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05511_ input4/X _11337_/Q _10213_/Q vssd1 vssd1 vccd1 vccd1 _11607_/D sky130_fd_sc_hd__mux2_1
X_06491_ _11871_/A _06485_/X _06490_/X _06576_/A vssd1 vssd1 vccd1 vccd1 _06491_/X
+ sky130_fd_sc_hd__a31o_1
X_05442_ _10506_/Q _09566_/D _09947_/B1 _10672_/Q vssd1 vssd1 vccd1 vccd1 _05442_/X
+ sky130_fd_sc_hd__a22o_1
X_08230_ _10137_/A _08230_/B _10087_/C vssd1 vssd1 vccd1 vccd1 _08325_/B sky130_fd_sc_hd__or3_4
XFILLER_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05373_ _05373_/A _05373_/B _05373_/C _05373_/D vssd1 vssd1 vccd1 vccd1 _05379_/A
+ sky130_fd_sc_hd__or4_4
X_08161_ _10106_/A1 _08162_/S _08160_/X _08843_/C1 vssd1 vssd1 vccd1 vccd1 _10906_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07112_ _07664_/A _07126_/B vssd1 vssd1 vccd1 vccd1 _07112_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08092_ _08092_/A _08655_/B vssd1 vssd1 vccd1 vccd1 _08092_/X sky130_fd_sc_hd__or2_4
XFILLER_107_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07043_ _09228_/A _07043_/B vssd1 vssd1 vccd1 vccd1 _07043_/X sky130_fd_sc_hd__or2_4
XFILLER_118_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08994_ _08994_/A _10180_/C _10137_/B vssd1 vssd1 vccd1 vccd1 _08994_/X sky130_fd_sc_hd__or3_4
XFILLER_141_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ _10787_/Q _07941_/Y _07944_/Y _08326_/B2 vssd1 vssd1 vccd1 vccd1 _10787_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07876_ _09182_/A0 _07890_/A2 _07875_/X _07932_/C1 vssd1 vssd1 vccd1 vccd1 _10756_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09615_ _09615_/A _09615_/B _09615_/C _09615_/D vssd1 vssd1 vccd1 vccd1 _09615_/X
+ sky130_fd_sc_hd__or4_2
X_06827_ _10375_/Q _07203_/A _06858_/B1 _10277_/Q vssd1 vssd1 vccd1 vccd1 _06827_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_70_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09546_ _05078_/A _09541_/Y _09545_/X _09833_/A vssd1 vssd1 vccd1 vccd1 _11625_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06758_ _10330_/Q _07111_/A _10009_/A _11716_/Q vssd1 vssd1 vccd1 vccd1 _06758_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_145_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05709_ _05709_/A _05709_/B _05709_/C _05709_/D vssd1 vssd1 vccd1 vccd1 _05716_/A
+ sky130_fd_sc_hd__or4_2
X_09477_ _09477_/A _09681_/B vssd1 vssd1 vccd1 vccd1 _09478_/C sky130_fd_sc_hd__nand2_1
XFILLER_12_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06689_ _10326_/Q _06856_/A2 _06686_/X _06688_/X _06997_/A vssd1 vssd1 vccd1 vccd1
+ _06689_/X sky130_fd_sc_hd__o2111a_1
XFILLER_145_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08428_ _11053_/Q _08424_/Y _08427_/Y _08440_/B2 vssd1 vssd1 vccd1 vccd1 _11053_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08359_ _07107_/A _08360_/S _08358_/X _09022_/C1 vssd1 vssd1 vccd1 vccd1 _11022_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ _11410_/CLK _11370_/D vssd1 vssd1 vccd1 vccd1 _11370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10321_ _10812_/CLK _10321_/D vssd1 vssd1 vccd1 vccd1 _10321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10252_ _11712_/CLK _10252_/D vssd1 vssd1 vccd1 vccd1 _10252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10183_ _10183_/A0 _11804_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _11804_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout260 _08529_/S vssd1 vssd1 vccd1 vccd1 _08537_/S sky130_fd_sc_hd__buf_6
Xfanout271 _08200_/X vssd1 vssd1 vccd1 vccd1 _08219_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_120_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout282 _07904_/X vssd1 vssd1 vccd1 vccd1 _09206_/B sky130_fd_sc_hd__buf_6
Xfanout293 _09200_/S vssd1 vssd1 vccd1 vccd1 _09193_/B sky130_fd_sc_hd__buf_8
XFILLER_75_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_104_wb_clk_i clkbuf_4_10__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11472_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11706_ _11706_/CLK _11706_/D vssd1 vssd1 vccd1 vccd1 _11706_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11637_ _11641_/CLK _11637_/D vssd1 vssd1 vccd1 vccd1 _11637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11568_ _11634_/CLK _11568_/D vssd1 vssd1 vccd1 vccd1 _11568_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10519_ _11474_/CLK _10519_/D vssd1 vssd1 vccd1 vccd1 _10519_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11499_ _11684_/CLK _11499_/D vssd1 vssd1 vccd1 vccd1 _11499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05991_ _10876_/Q _06468_/B _06152_/B _10613_/Q _07083_/B vssd1 vssd1 vccd1 vccd1
+ _05991_/X sky130_fd_sc_hd__o221a_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07730_ _10666_/Q _07750_/B vssd1 vssd1 vccd1 vccd1 _07730_/X sky130_fd_sc_hd__or2_1
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07661_ _10624_/Q _07663_/S _07246_/S _07316_/B vssd1 vssd1 vccd1 vccd1 _10624_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09400_ _10105_/A1 _11566_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _11566_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06612_ _06606_/X _06611_/X _11872_/A vssd1 vssd1 vccd1 vccd1 _06612_/X sky130_fd_sc_hd__a21o_1
XFILLER_129_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07592_ _10056_/A _07592_/B vssd1 vssd1 vccd1 vccd1 _10579_/D sky130_fd_sc_hd__or2_1
XFILLER_52_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09331_ _11520_/Q _09343_/B vssd1 vssd1 vccd1 vccd1 _09331_/X sky130_fd_sc_hd__or2_1
XFILLER_94_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06543_ _11149_/Q _07692_/A _06629_/B1 _11100_/Q _07690_/B vssd1 vssd1 vccd1 vccd1
+ _06543_/X sky130_fd_sc_hd__o221a_2
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09262_ _10150_/A1 _09266_/B _08761_/A vssd1 vssd1 vccd1 vccd1 _09262_/X sky130_fd_sc_hd__a21o_1
X_06474_ _06461_/X _06462_/X _06473_/X _06619_/A1 vssd1 vssd1 vccd1 vccd1 _06474_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08213_ _09323_/A0 _10941_/Q _08225_/S vssd1 vssd1 vccd1 vccd1 _08214_/B sky130_fd_sc_hd__mux2_1
X_05425_ _11149_/Q _11148_/Q _09680_/C vssd1 vssd1 vccd1 vccd1 _05428_/B sky130_fd_sc_hd__mux2_1
X_09193_ _09193_/A _09193_/B vssd1 vssd1 vccd1 vccd1 _09193_/Y sky130_fd_sc_hd__nand2_4
XFILLER_147_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05356_ _05356_/A _05356_/B _05356_/C _05356_/D vssd1 vssd1 vccd1 vccd1 _05357_/B
+ sky130_fd_sc_hd__or4_4
X_08144_ _10898_/Q _08637_/C vssd1 vssd1 vccd1 vccd1 _08144_/X sky130_fd_sc_hd__or2_1
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05287_ _05085_/Y _11174_/Q _10899_/Q _09680_/B vssd1 vssd1 vccd1 vccd1 _05291_/C
+ sky130_fd_sc_hd__a22o_1
X_08075_ _10863_/Q _08085_/B vssd1 vssd1 vccd1 vccd1 _08075_/X sky130_fd_sc_hd__or2_1
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07026_ _09229_/A _07026_/B vssd1 vssd1 vccd1 vccd1 _07026_/X sky130_fd_sc_hd__and2_2
XFILLER_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08977_ _11341_/Q _08989_/B vssd1 vssd1 vccd1 vccd1 _08977_/X sky130_fd_sc_hd__or2_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11262_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07928_ _07928_/A _07928_/B vssd1 vssd1 vccd1 vccd1 _10781_/D sky130_fd_sc_hd__or2_1
XFILLER_57_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07859_ _10748_/Q _07883_/B vssd1 vssd1 vccd1 vccd1 _07859_/X sky130_fd_sc_hd__or2_1
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10870_ _11633_/CLK _10870_/D vssd1 vssd1 vccd1 vccd1 _10870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09529_/A _09529_/B _09529_/C vssd1 vssd1 vccd1 vccd1 _11619_/D sky130_fd_sc_hd__and3_1
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11422_ _11428_/CLK _11422_/D vssd1 vssd1 vccd1 vccd1 _11422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11353_ _11366_/CLK _11353_/D vssd1 vssd1 vccd1 vccd1 _11353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10304_ _11768_/CLK _10304_/D vssd1 vssd1 vccd1 vccd1 _10304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11284_ _11284_/CLK _11284_/D vssd1 vssd1 vccd1 vccd1 _11284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10235_ _11657_/CLK _10235_/D vssd1 vssd1 vccd1 vccd1 _10235_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_105_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1000 input82/X vssd1 vssd1 vccd1 vccd1 _06357_/C1 sky130_fd_sc_hd__clkbuf_16
XFILLER_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1011 _10178_/A1 vssd1 vssd1 vccd1 vccd1 _09101_/A1 sky130_fd_sc_hd__buf_6
XFILLER_120_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1022 _10177_/A1 vssd1 vssd1 vccd1 vccd1 _09214_/A sky130_fd_sc_hd__buf_6
XFILLER_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10166_ _10166_/A1 _10176_/B _10166_/B1 vssd1 vssd1 vccd1 vccd1 _10166_/X sky130_fd_sc_hd__a21o_1
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1033 input114/X vssd1 vssd1 vccd1 vccd1 _07015_/A sky130_fd_sc_hd__buf_6
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1044 _08919_/A1 vssd1 vssd1 vccd1 vccd1 _10019_/A0 sky130_fd_sc_hd__buf_12
Xfanout1055 _10184_/A0 vssd1 vssd1 vccd1 vccd1 _09395_/A0 sky130_fd_sc_hd__clkbuf_8
Xfanout1066 _10142_/A1 vssd1 vssd1 vccd1 vccd1 _07007_/A sky130_fd_sc_hd__buf_12
Xfanout1077 input101/X vssd1 vssd1 vccd1 vccd1 _07034_/A sky130_fd_sc_hd__buf_6
XFILLER_43_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10097_ _11750_/Q _10087_/X _10096_/X vssd1 vssd1 vccd1 vccd1 _11750_/D sky130_fd_sc_hd__a21o_1
XFILLER_78_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10999_ _11763_/CLK _10999_/D vssd1 vssd1 vccd1 vccd1 _10999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05210_ _10906_/Q _10905_/Q _06945_/B vssd1 vssd1 vccd1 vccd1 _05213_/B sky130_fd_sc_hd__mux2_1
X_06190_ _11465_/Q _07152_/A vssd1 vssd1 vccd1 vccd1 _06190_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_72_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11497_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_156_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05141_ _10634_/Q _10633_/Q _05418_/S vssd1 vssd1 vccd1 vccd1 _05145_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05072_ _09497_/A vssd1 vssd1 vccd1 vccd1 _05072_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08900_ _11309_/Q _07100_/X _08901_/S vssd1 vssd1 vccd1 vccd1 _11309_/D sky130_fd_sc_hd__mux2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _09880_/A _09880_/B _09880_/C _09880_/D vssd1 vssd1 vccd1 vccd1 _09888_/B
+ sky130_fd_sc_hd__or4_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08969_/A1 _08832_/S _08830_/X _08831_/C1 vssd1 vssd1 vccd1 vccd1 _11273_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _11238_/Q _08762_/B vssd1 vssd1 vccd1 vccd1 _08762_/X sky130_fd_sc_hd__or2_1
XFILLER_22_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05974_ _10656_/Q _07455_/A vssd1 vssd1 vccd1 vccd1 _05974_/X sky130_fd_sc_hd__or2_1
XFILLER_61_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07713_ _10017_/A0 _07755_/A2 _07712_/X _07868_/C1 vssd1 vssd1 vccd1 vccd1 _10657_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_tms1x00_1109 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1109/HI io_out[1] sky130_fd_sc_hd__conb_1
X_08693_ _11201_/Q _08705_/B vssd1 vssd1 vccd1 vccd1 _08693_/X sky130_fd_sc_hd__or2_1
XFILLER_93_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07644_ _08193_/A _08197_/S vssd1 vssd1 vccd1 vccd1 _07644_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07575_ _07028_/A _10571_/Q _07593_/S vssd1 vssd1 vccd1 vccd1 _07576_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09314_ _09314_/A _10108_/B _10119_/C vssd1 vssd1 vccd1 vccd1 _09324_/S sky130_fd_sc_hd__or3_4
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06526_ _10356_/Q _08649_/A _06523_/X _06525_/X vssd1 vssd1 vccd1 vccd1 _06526_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_55_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09245_ _11475_/Q _09226_/Y _09229_/Y _07451_/X vssd1 vssd1 vccd1 vccd1 _11475_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06457_ _10829_/Q _07994_/A _06628_/B1 _11274_/Q vssd1 vssd1 vccd1 vccd1 _06457_/X
+ sky130_fd_sc_hd__o22a_1
X_05408_ _11282_/Q _11281_/Q _05419_/S vssd1 vssd1 vccd1 vccd1 _05411_/B sky130_fd_sc_hd__mux2_1
X_09176_ _09193_/A _09187_/S vssd1 vssd1 vccd1 vccd1 _09176_/Y sky130_fd_sc_hd__nand2_2
X_06388_ _10894_/Q _08123_/A vssd1 vssd1 vccd1 vccd1 _06388_/X sky130_fd_sc_hd__or2_1
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08127_ _08590_/A _08127_/B vssd1 vssd1 vccd1 vccd1 _10889_/D sky130_fd_sc_hd__or2_1
X_05339_ _11088_/Q _11087_/Q _05427_/S vssd1 vssd1 vccd1 vccd1 _05340_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08058_ _10190_/A0 _08427_/B _08057_/X _08345_/C1 vssd1 vssd1 vccd1 vccd1 _10854_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07009_ _10267_/Q _07008_/X _07038_/S vssd1 vssd1 vccd1 vccd1 _10267_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10020_ _10020_/A _10020_/B vssd1 vssd1 vccd1 vccd1 _11700_/D sky130_fd_sc_hd__or2_1
Xinput103 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 input103/X sky130_fd_sc_hd__clkbuf_8
Xinput114 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 input114/X sky130_fd_sc_hd__buf_6
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ _11220_/CLK _10922_/D vssd1 vssd1 vccd1 vccd1 _10922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10853_ _11023_/CLK _10853_/D vssd1 vssd1 vccd1 vccd1 _10853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10784_ _11439_/CLK _10784_/D vssd1 vssd1 vccd1 vccd1 _10784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11405_ _11411_/CLK _11405_/D vssd1 vssd1 vccd1 vccd1 _11405_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_153_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11336_ _11675_/CLK _11336_/D vssd1 vssd1 vccd1 vccd1 _11336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11267_ _11779_/CLK _11267_/D vssd1 vssd1 vccd1 vccd1 _11267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10218_ _10765_/CLK _10218_/D vssd1 vssd1 vccd1 vccd1 _10218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11198_ _11319_/CLK _11198_/D vssd1 vssd1 vccd1 vccd1 _11198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10149_ _10149_/A1 _10137_/X _10148_/X _10153_/C1 vssd1 vssd1 vccd1 vccd1 _11787_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05690_ _11157_/Q _05609_/Y _05615_/Y _11165_/Q _05689_/X vssd1 vssd1 vccd1 vccd1
+ _05691_/C sky130_fd_sc_hd__a221o_1
XFILLER_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07360_ _08440_/B2 _10451_/Q _07363_/S vssd1 vssd1 vccd1 vccd1 _10451_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06311_ _11041_/Q _08383_/A _06363_/A2 _10963_/Q vssd1 vssd1 vccd1 vccd1 _06311_/X
+ sky130_fd_sc_hd__o22a_1
X_07291_ _07036_/A _10414_/Q _09184_/S vssd1 vssd1 vccd1 vccd1 _07292_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09030_ _10150_/A1 _09016_/X _09029_/X _09036_/C1 vssd1 vssd1 vccd1 vccd1 _11365_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06242_ _11434_/Q _06804_/B _07455_/A _10660_/Q vssd1 vssd1 vccd1 vccd1 _06242_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06173_ _11345_/Q _08972_/A _06716_/B1 _11408_/Q vssd1 vssd1 vccd1 vccd1 _06173_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05124_ _05124_/A _05124_/B vssd1 vssd1 vccd1 vccd1 _05124_/Y sky130_fd_sc_hd__nor2_4
X_09932_ _11659_/Q _09770_/S _09929_/X _09931_/X vssd1 vssd1 vccd1 vccd1 _11659_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout804 _06351_/A2 vssd1 vssd1 vccd1 vccd1 _10072_/A sky130_fd_sc_hd__buf_4
Xfanout815 _06166_/A2 vssd1 vssd1 vccd1 vccd1 _06412_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout826 _06238_/A2 vssd1 vssd1 vccd1 vccd1 _06470_/A2 sky130_fd_sc_hd__buf_4
Xfanout837 _06803_/A2 vssd1 vssd1 vccd1 vccd1 _06872_/A2 sky130_fd_sc_hd__buf_6
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _10706_/Q _09573_/A _09567_/B _11445_/Q vssd1 vssd1 vccd1 vccd1 _09863_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout848 _10086_/A vssd1 vssd1 vccd1 vccd1 _06648_/A2 sky130_fd_sc_hd__clkbuf_16
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout859 _06230_/A2 vssd1 vssd1 vccd1 vccd1 _06540_/A2 sky130_fd_sc_hd__buf_6
X_08814_ _11264_/Q _08820_/S _07630_/Y _07098_/B vssd1 vssd1 vccd1 vccd1 _11264_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09794_ _11651_/Q _08950_/B _09793_/X _09478_/A vssd1 vssd1 vccd1 vccd1 _11651_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08745_ _08745_/A _08745_/B vssd1 vssd1 vccd1 vccd1 _11229_/D sky130_fd_sc_hd__or2_1
XFILLER_100_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05957_ _11392_/Q _06716_/A2 _06717_/B1 _11342_/Q vssd1 vssd1 vccd1 vccd1 _05957_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_6_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _07018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _08793_/A _08676_/B vssd1 vssd1 vccd1 vccd1 _11192_/D sky130_fd_sc_hd__or2_1
X_05888_ _11748_/Q _10087_/A _10137_/A _11784_/Q _06349_/C1 vssd1 vssd1 vccd1 vccd1
+ _05888_/X sky130_fd_sc_hd__o221a_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _07108_/X _10599_/Q _07628_/S vssd1 vssd1 vccd1 vccd1 _10599_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07558_ _08684_/A _07558_/B vssd1 vssd1 vccd1 vccd1 _10562_/D sky130_fd_sc_hd__or2_1
X_06509_ _10884_/Q _06468_/B _06508_/X _06642_/C1 vssd1 vssd1 vccd1 vccd1 _06509_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07489_ _07105_/X _10525_/Q _07490_/S vssd1 vssd1 vccd1 vccd1 _10525_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09228_ _09228_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09159_ _11424_/Q _09171_/B vssd1 vssd1 vccd1 vccd1 _09159_/X sky130_fd_sc_hd__or2_1
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11121_ _11291_/CLK _11121_/D vssd1 vssd1 vccd1 vccd1 _11121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11052_ _11572_/CLK _11052_/D vssd1 vssd1 vccd1 vccd1 _11052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10003_ _10113_/A0 _11690_/Q _10008_/S vssd1 vssd1 vccd1 vccd1 _11690_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10905_ _11235_/CLK _10905_/D vssd1 vssd1 vccd1 vccd1 _10905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10836_ _11243_/CLK _10836_/D vssd1 vssd1 vccd1 vccd1 _10836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10767_ _11462_/CLK _10767_/D vssd1 vssd1 vccd1 vccd1 _10767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10698_ _11622_/CLK _10698_/D vssd1 vssd1 vccd1 vccd1 _10698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11319_ _11319_/CLK _11319_/D vssd1 vssd1 vccd1 vccd1 _11319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06860_ _10631_/Q _06860_/A2 _06856_/X _06859_/X vssd1 vssd1 vccd1 vccd1 _06860_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05811_ _10645_/Q _07692_/A _05809_/X _05810_/X vssd1 vssd1 vccd1 vccd1 _05811_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06791_ _10715_/Q _07778_/A _06805_/B1 _10550_/Q vssd1 vssd1 vccd1 vccd1 _06791_/X
+ sky130_fd_sc_hd__o22a_1
X_08530_ _08783_/A _08530_/B vssd1 vssd1 vccd1 vccd1 _11114_/D sky130_fd_sc_hd__or2_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05742_ _05745_/A _05749_/A _05751_/B vssd1 vssd1 vccd1 vccd1 _05742_/Y sky130_fd_sc_hd__nor3_4
XFILLER_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08461_ _11081_/Q _10128_/A0 _08467_/S vssd1 vssd1 vccd1 vccd1 _08462_/B sky130_fd_sc_hd__mux2_1
X_05673_ _11205_/Q _05579_/Y _05597_/Y _11196_/Q _05669_/X vssd1 vssd1 vccd1 vccd1
+ _05680_/A sky130_fd_sc_hd__a221o_1
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07412_ _10026_/A _07412_/B vssd1 vssd1 vccd1 vccd1 _10482_/D sky130_fd_sc_hd__or2_1
XFILLER_56_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08392_ _09141_/A1 _11037_/Q _08414_/S vssd1 vssd1 vccd1 vccd1 _08393_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07343_ _10439_/Q _07337_/X _07846_/S _07229_/B vssd1 vssd1 vccd1 vccd1 _10439_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07274_ _08883_/A1 _07277_/S _07273_/X _07894_/C1 vssd1 vssd1 vccd1 vccd1 _10405_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09013_ _11358_/Q _09013_/B vssd1 vssd1 vccd1 vccd1 _09013_/X sky130_fd_sc_hd__or2_1
X_06225_ _11730_/Q _10061_/A _09347_/A _11535_/Q vssd1 vssd1 vccd1 vccd1 _06225_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06156_ _10915_/Q _06591_/A2 _06155_/X _11869_/A vssd1 vssd1 vccd1 vccd1 _06156_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05107_ _05107_/A _05107_/B _05107_/C _05107_/D vssd1 vssd1 vccd1 vccd1 _05113_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06087_ _11681_/Q _09977_/A _06083_/X _06086_/X vssd1 vssd1 vccd1 vccd1 _06093_/B
+ sky130_fd_sc_hd__o211a_1
Xfanout601 _05774_/Y vssd1 vssd1 vccd1 vccd1 _06743_/B sky130_fd_sc_hd__buf_4
Xfanout612 _07300_/A vssd1 vssd1 vccd1 vccd1 _06228_/A2 sky130_fd_sc_hd__buf_4
XFILLER_132_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09915_ _10485_/Q _09947_/A2 _09568_/C _10357_/Q vssd1 vssd1 vccd1 vccd1 _09915_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout623 _06696_/A2 vssd1 vssd1 vccd1 vccd1 _08383_/A sky130_fd_sc_hd__buf_4
XFILLER_63_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout634 _09529_/A vssd1 vssd1 vccd1 vccd1 _09825_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout645 _05076_/Y vssd1 vssd1 vccd1 vccd1 _05616_/A1 sky130_fd_sc_hd__buf_6
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout656 _11653_/Q vssd1 vssd1 vccd1 vccd1 _09515_/C sky130_fd_sc_hd__buf_4
XFILLER_115_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09846_ _10770_/Q _09875_/A2 _09872_/A2 _10785_/Q vssd1 vssd1 vccd1 vccd1 _09846_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout667 _09430_/B vssd1 vssd1 vccd1 vccd1 _05399_/S sky130_fd_sc_hd__buf_8
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout678 _05430_/S vssd1 vssd1 vccd1 vccd1 _05398_/S sky130_fd_sc_hd__buf_4
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 _05326_/S vssd1 vssd1 vccd1 vccd1 _05414_/S sky130_fd_sc_hd__buf_6
XFILLER_101_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _09404_/Y _09775_/X _09776_/Y _09681_/B vssd1 vssd1 vccd1 vccd1 _09777_/X
+ sky130_fd_sc_hd__a31o_1
X_06989_ _10262_/Q _06995_/B vssd1 vssd1 vccd1 vccd1 _06989_/X sky130_fd_sc_hd__or2_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _07007_/A _11221_/Q _08742_/S vssd1 vssd1 vccd1 vccd1 _08729_/B sky130_fd_sc_hd__mux2_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _11185_/Q _07104_/A _08663_/S vssd1 vssd1 vccd1 vccd1 _08660_/B sky130_fd_sc_hd__mux2_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11758_/CLK _11670_/D vssd1 vssd1 vccd1 vccd1 _11670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10621_ _11702_/CLK _10621_/D vssd1 vssd1 vccd1 vccd1 _10621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ _10769_/CLK _10552_/D vssd1 vssd1 vccd1 vccd1 _10552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10483_ _11710_/CLK _10483_/D vssd1 vssd1 vccd1 vccd1 _10483_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_129_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10812_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11104_ _11393_/CLK _11104_/D vssd1 vssd1 vccd1 vccd1 _11104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11035_ _11683_/CLK _11035_/D vssd1 vssd1 vccd1 vccd1 _11035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11868_ _11868_/A vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__buf_2
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10819_ _10932_/CLK _10819_/D vssd1 vssd1 vccd1 vccd1 _10819_/Q sky130_fd_sc_hd__dfxtp_1
X_11799_ _11801_/CLK _11799_/D vssd1 vssd1 vccd1 vccd1 _11799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06010_ _10950_/Q _06504_/B1 _06006_/X _06009_/X vssd1 vssd1 vccd1 vccd1 _06010_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput204 _05508_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_4
XFILLER_154_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07961_ _07040_/X _10803_/Q _07961_/S vssd1 vssd1 vccd1 vccd1 _10803_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _11637_/Q _11641_/Q _09702_/S vssd1 vssd1 vccd1 vccd1 _09701_/B sky130_fd_sc_hd__mux2_1
X_06912_ _10197_/Q _06922_/B vssd1 vssd1 vccd1 vccd1 _06912_/X sky130_fd_sc_hd__or2_1
X_07892_ _07933_/A0 _07966_/S _07891_/X _07902_/C1 vssd1 vssd1 vccd1 vccd1 _10764_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09631_ _10734_/Q _09572_/B _09572_/C _10735_/Q _09627_/X vssd1 vssd1 vccd1 vccd1
+ _09633_/C sky130_fd_sc_hd__a221o_1
X_06843_ _10767_/Q _07854_/A _06875_/B1 _10506_/Q vssd1 vssd1 vccd1 vccd1 _06843_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09562_ _11659_/Q _11644_/Q vssd1 vssd1 vccd1 vccd1 _09564_/A sky130_fd_sc_hd__and2_2
X_06774_ _10360_/Q _06803_/A2 _06773_/X _06849_/C1 vssd1 vssd1 vccd1 vccd1 _06774_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08513_ _11106_/Q _08545_/B vssd1 vssd1 vccd1 vccd1 _08513_/X sky130_fd_sc_hd__or2_1
X_05725_ _10960_/Q _05609_/Y _05627_/Y _10955_/Q _05724_/X vssd1 vssd1 vccd1 vccd1
+ _05728_/C sky130_fd_sc_hd__a221o_2
X_09493_ _11609_/Q _09490_/Y _09492_/X _09529_/A vssd1 vssd1 vccd1 vccd1 _11609_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08444_ _11065_/Q _08436_/Y _08439_/Y _07316_/X vssd1 vssd1 vccd1 vccd1 _11065_/D
+ sky130_fd_sc_hd__a22o_1
X_05656_ _11289_/Q _05603_/Y _05653_/X _05655_/X vssd1 vssd1 vccd1 vccd1 _05656_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_23_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08375_ _10150_/A1 _08439_/B _08374_/X _08662_/C1 vssd1 vssd1 vccd1 vccd1 _11029_/D
+ sky130_fd_sc_hd__o211a_1
X_05587_ _05629_/A2 _10201_/Q _10195_/Q _05629_/B1 vssd1 vssd1 vccd1 vccd1 _05587_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07326_ _08439_/A _08162_/S vssd1 vssd1 vccd1 vccd1 _07326_/Y sky130_fd_sc_hd__nand2_4
XFILLER_104_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07257_ _10013_/A0 _10397_/Q _09187_/S vssd1 vssd1 vccd1 vccd1 _07258_/B sky130_fd_sc_hd__mux2_1
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06208_ _07082_/A _06206_/X _06207_/X _06576_/A vssd1 vssd1 vccd1 vccd1 _06208_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07188_ _07187_/X _10355_/Q _07188_/S vssd1 vssd1 vccd1 vccd1 _10355_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06139_ _10420_/Q _06318_/A2 _06538_/A2 _11028_/Q _06138_/X vssd1 vssd1 vccd1 vccd1
+ _06139_/X sky130_fd_sc_hd__o221a_1
XFILLER_79_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout420 _05313_/Y vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_63_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout431 _05259_/Y vssd1 vssd1 vccd1 vccd1 _09883_/B1 sky130_fd_sc_hd__buf_4
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout442 _05190_/Y vssd1 vssd1 vccd1 vccd1 _09568_/B sky130_fd_sc_hd__buf_8
Xfanout453 _05135_/Y vssd1 vssd1 vccd1 vccd1 _09879_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout464 _08345_/C1 vssd1 vssd1 vccd1 vccd1 _08351_/C1 sky130_fd_sc_hd__buf_4
XFILLER_101_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout475 _10155_/C1 vssd1 vssd1 vccd1 vccd1 _09267_/C1 sky130_fd_sc_hd__buf_4
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout486 _07884_/C1 vssd1 vssd1 vccd1 vccd1 _07894_/C1 sky130_fd_sc_hd__buf_4
XFILLER_101_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout497 _09168_/C1 vssd1 vssd1 vccd1 vccd1 _10175_/C1 sky130_fd_sc_hd__buf_4
XFILLER_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09829_ _09824_/S _09827_/Y _09828_/Y vssd1 vssd1 vccd1 vccd1 _11656_/D sky130_fd_sc_hd__a21oi_1
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11722_ _11722_/CLK _11722_/D vssd1 vssd1 vccd1 vccd1 _11722_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11663_/CLK _11653_/D vssd1 vssd1 vccd1 vccd1 _11653_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ _11262_/CLK _10604_/D vssd1 vssd1 vccd1 vccd1 _10604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ _11584_/CLK _11584_/D vssd1 vssd1 vccd1 vccd1 _11584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10535_ _10805_/CLK _10535_/D vssd1 vssd1 vccd1 vccd1 _10535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10466_ _10981_/CLK _10466_/D vssd1 vssd1 vccd1 vccd1 _10466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10397_ _10804_/CLK _10397_/D vssd1 vssd1 vccd1 vccd1 _10397_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_6_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_97_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _10805_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11018_ _11023_/CLK _11018_/D vssd1 vssd1 vccd1 vccd1 _11018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_26_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11632_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05510_ input3/X _11336_/Q _10213_/Q vssd1 vssd1 vccd1 vccd1 _11606_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06490_ _11163_/Q _06649_/A2 _06486_/X _06489_/X vssd1 vssd1 vccd1 vccd1 _06490_/X
+ sky130_fd_sc_hd__a211o_4
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05441_ _10505_/Q _09566_/B _09568_/D _10655_/Q _05440_/X vssd1 vssd1 vccd1 vccd1
+ _05451_/B sky130_fd_sc_hd__a221o_1
XFILLER_18_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08160_ _10906_/Q _08164_/B vssd1 vssd1 vccd1 vccd1 _08160_/X sky130_fd_sc_hd__or2_1
XFILLER_18_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05372_ _10825_/Q _10824_/Q _05372_/S vssd1 vssd1 vccd1 vccd1 _05373_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07111_ _07111_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _07111_/X sky130_fd_sc_hd__or2_4
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08091_ _10871_/Q _08655_/B _08091_/C vssd1 vssd1 vccd1 vccd1 _08091_/X sky130_fd_sc_hd__or3_1
XFILLER_88_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07042_ _07042_/A _07205_/A vssd1 vssd1 vccd1 vccd1 _07043_/B sky130_fd_sc_hd__and2_2
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08993_ _10136_/A _09015_/B _10158_/B vssd1 vssd1 vccd1 vccd1 _09013_/B sky130_fd_sc_hd__and3_4
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07944_ _08439_/A _08083_/S vssd1 vssd1 vccd1 vccd1 _07944_/Y sky130_fd_sc_hd__nand2_2
XFILLER_60_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07875_ _10756_/Q _07893_/B vssd1 vssd1 vccd1 vccd1 _07875_/X sky130_fd_sc_hd__or2_1
XFILLER_56_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06826_ _11333_/Q _06704_/B _06825_/X vssd1 vssd1 vccd1 vccd1 _10247_/D sky130_fd_sc_hd__a21o_1
X_09614_ _10620_/Q _09566_/B _09573_/B _10624_/Q _09601_/X vssd1 vssd1 vccd1 vccd1
+ _09615_/D sky130_fd_sc_hd__a221o_2
XFILLER_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09545_ _11663_/Q _09538_/X _09542_/X vssd1 vssd1 vccd1 vccd1 _09545_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06757_ _10373_/Q _07203_/A _06858_/B1 _10276_/Q vssd1 vssd1 vccd1 vccd1 _06757_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05708_ _11035_/Q _05531_/Y _05555_/Y _11044_/Q vssd1 vssd1 vccd1 vccd1 _05709_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_145_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09476_ _09680_/B _09407_/B _09475_/Y _09478_/A vssd1 vssd1 vccd1 vccd1 _11601_/D
+ sky130_fd_sc_hd__o211a_1
X_06688_ _10292_/Q _06873_/A2 _06858_/B1 _10274_/Q _06687_/X vssd1 vssd1 vccd1 vccd1
+ _06688_/X sky130_fd_sc_hd__o221a_1
XFILLER_58_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08427_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08427_/Y sky130_fd_sc_hd__nand2_2
XFILLER_145_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05639_ _11315_/Q _05531_/Y _05567_/Y _11316_/Q vssd1 vssd1 vccd1 vccd1 _05639_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08358_ _11022_/Q _08362_/B vssd1 vssd1 vccd1 vccd1 _08358_/X sky130_fd_sc_hd__or2_1
XFILLER_149_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07309_ _07309_/A _07617_/B vssd1 vssd1 vccd1 vccd1 _07309_/X sky130_fd_sc_hd__or2_4
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08289_ _10975_/Q _07088_/X _08298_/S vssd1 vssd1 vccd1 vccd1 _10975_/D sky130_fd_sc_hd__mux2_1
XFILLER_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10320_ _10812_/CLK _10320_/D vssd1 vssd1 vccd1 vccd1 _10320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _11712_/CLK _10251_/D vssd1 vssd1 vccd1 vccd1 _10251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10182_ _10182_/A0 _11803_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _11803_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout250 _08855_/X vssd1 vssd1 vccd1 vccd1 _08874_/S sky130_fd_sc_hd__buf_6
XFILLER_59_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout261 _08506_/X vssd1 vssd1 vccd1 vccd1 _08529_/S sky130_fd_sc_hd__buf_8
Xfanout272 _08166_/X vssd1 vssd1 vccd1 vccd1 _08181_/S sky130_fd_sc_hd__buf_6
Xfanout283 _07890_/A2 vssd1 vssd1 vccd1 vccd1 _07966_/S sky130_fd_sc_hd__buf_6
XFILLER_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout294 _09200_/S vssd1 vssd1 vccd1 vccd1 _07817_/S sky130_fd_sc_hd__buf_8
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11705_ _11720_/CLK _11705_/D vssd1 vssd1 vccd1 vccd1 _11705_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11636_ _11641_/CLK _11636_/D vssd1 vssd1 vccd1 vccd1 _11636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11567_ _11675_/CLK _11567_/D vssd1 vssd1 vccd1 vccd1 _11567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10518_ _11474_/CLK _10518_/D vssd1 vssd1 vccd1 vccd1 _10518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11498_ _11801_/CLK _11498_/D vssd1 vssd1 vccd1 vccd1 _11498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10449_ _11133_/CLK _10449_/D vssd1 vssd1 vccd1 vccd1 _10449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05990_ _10458_/Q _06308_/A2 _07111_/A _10811_/Q vssd1 vssd1 vccd1 vccd1 _05990_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07660_ _10623_/Q _07663_/S _07246_/S _07314_/B vssd1 vssd1 vccd1 vccd1 _10623_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_66_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06611_ _11709_/Q _08560_/A _06607_/X _06610_/X vssd1 vssd1 vccd1 vccd1 _06611_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_19_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07591_ _07143_/A _10579_/Q _07591_/S vssd1 vssd1 vccd1 vccd1 _07592_/B sky130_fd_sc_hd__mux2_1
XFILLER_81_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ _10162_/A1 _09326_/X _09329_/X _09993_/C1 vssd1 vssd1 vccd1 vccd1 _11519_/D
+ sky130_fd_sc_hd__o211a_1
X_06542_ _10831_/Q _07994_/A _06628_/B1 _11276_/Q vssd1 vssd1 vccd1 vccd1 _06542_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09261_ _11483_/Q _09249_/X _09260_/X vssd1 vssd1 vccd1 vccd1 _11483_/D sky130_fd_sc_hd__a21o_1
XFILLER_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06473_ _06469_/X _06472_/X _07083_/A _06467_/X vssd1 vssd1 vccd1 vccd1 _06473_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08212_ _08492_/A _08212_/B vssd1 vssd1 vccd1 vccd1 _10940_/D sky130_fd_sc_hd__or2_1
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05424_ _10647_/Q _11147_/Q _11596_/Q vssd1 vssd1 vccd1 vccd1 _05428_/A sky130_fd_sc_hd__mux2_1
X_09192_ _09192_/A _09192_/B vssd1 vssd1 vccd1 vccd1 _09192_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08143_ _08835_/A _08143_/B vssd1 vssd1 vccd1 vccd1 _10897_/D sky130_fd_sc_hd__or2_1
X_05355_ _11136_/Q _11135_/Q _05391_/S vssd1 vssd1 vccd1 vccd1 _05356_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08074_ _10015_/A0 _08083_/S _08073_/X _08753_/C1 vssd1 vssd1 vccd1 vccd1 _10862_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05286_ _06941_/A _10900_/Q _10893_/Q _05377_/S vssd1 vssd1 vccd1 vccd1 _05291_/B
+ sky130_fd_sc_hd__a22o_2
X_07025_ _07025_/A _07928_/A vssd1 vssd1 vccd1 vccd1 _07026_/B sky130_fd_sc_hd__or2_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08976_ _11340_/Q _08972_/X _08975_/X vssd1 vssd1 vccd1 vccd1 _11340_/D sky130_fd_sc_hd__a21o_1
XFILLER_64_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07927_ _07031_/A _10781_/Q _09221_/C vssd1 vssd1 vccd1 vccd1 _07928_/B sky130_fd_sc_hd__mux2_1
XFILLER_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07858_ _10013_/A0 _07871_/S _07857_/X _07868_/C1 vssd1 vssd1 vccd1 vccd1 _10747_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06809_ _06804_/X _06805_/X _06808_/X _06803_/X vssd1 vssd1 vccd1 vccd1 _06809_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07789_ _10019_/A0 _10702_/Q _07817_/S vssd1 vssd1 vccd1 vccd1 _07790_/B sky130_fd_sc_hd__mux2_1
XFILLER_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _09528_/A _09528_/B _09500_/C vssd1 vssd1 vccd1 vccd1 _09529_/C sky130_fd_sc_hd__or3b_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09441_/A input13/X _09441_/B vssd1 vssd1 vccd1 vccd1 _09459_/X sky130_fd_sc_hd__o21a_1
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _11792_/CLK _11421_/D vssd1 vssd1 vccd1 vccd1 _11421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11352_ _11366_/CLK _11352_/D vssd1 vssd1 vccd1 vccd1 _11352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10303_ _11776_/CLK _10303_/D vssd1 vssd1 vccd1 vccd1 _10303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11283_ _11527_/CLK _11283_/D vssd1 vssd1 vccd1 vccd1 _11283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10234_ _11665_/CLK _10234_/D vssd1 vssd1 vccd1 vccd1 _10234_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_152_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1001 _11868_/A vssd1 vssd1 vccd1 vccd1 _05751_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_79_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1012 _09129_/A1 vssd1 vssd1 vccd1 vccd1 _10178_/A1 sky130_fd_sc_hd__clkbuf_16
X_10165_ _10165_/A1 _10159_/X _10164_/X _10177_/C1 vssd1 vssd1 vccd1 vccd1 _11794_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout1023 input116/X vssd1 vssd1 vccd1 vccd1 _10177_/A1 sky130_fd_sc_hd__buf_12
Xfanout1034 _09124_/A1 vssd1 vssd1 vccd1 vccd1 _09285_/A1 sky130_fd_sc_hd__buf_6
Xfanout1045 input113/X vssd1 vssd1 vccd1 vccd1 _08919_/A1 sky130_fd_sc_hd__buf_12
XFILLER_43_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1056 _10184_/A0 vssd1 vssd1 vccd1 vccd1 _09256_/A1 sky130_fd_sc_hd__buf_6
XFILLER_82_1291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10096_ _10185_/A0 _10104_/B _10156_/B1 vssd1 vssd1 vccd1 vccd1 _10096_/X sky130_fd_sc_hd__a21o_1
Xfanout1067 _10165_/A1 vssd1 vssd1 vccd1 vccd1 _09364_/A1 sky130_fd_sc_hd__buf_6
Xfanout1078 input100/X vssd1 vssd1 vccd1 vccd1 _10047_/A1 sky130_fd_sc_hd__buf_6
XFILLER_47_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10998_ _11735_/CLK _10998_/D vssd1 vssd1 vccd1 vccd1 _10998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11619_ _11622_/CLK _11619_/D vssd1 vssd1 vccd1 vccd1 _11619_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05140_ _05140_/A _05140_/B _05140_/C _05140_/D vssd1 vssd1 vccd1 vccd1 _05146_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_41_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11811_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08830_ _11273_/Q _08840_/B vssd1 vssd1 vccd1 vccd1 _08830_/X sky130_fd_sc_hd__or2_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08761_/A _08761_/B vssd1 vssd1 vccd1 vccd1 _11237_/D sky130_fd_sc_hd__or2_1
X_05973_ _06189_/A1 _05967_/X _05972_/X _08243_/A _05962_/X vssd1 vssd1 vccd1 vccd1
+ _05973_/X sky130_fd_sc_hd__o311a_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07712_ _10657_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07712_/X sky130_fd_sc_hd__or2_1
XFILLER_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08692_ _08771_/A _08692_/B vssd1 vssd1 vccd1 vccd1 _11200_/D sky130_fd_sc_hd__or2_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07643_ _09976_/A _08649_/B _07643_/C vssd1 vssd1 vccd1 vccd1 _07645_/B sky130_fd_sc_hd__and3_2
XFILLER_54_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07574_ _07930_/A _07574_/B vssd1 vssd1 vccd1 vccd1 _10570_/D sky130_fd_sc_hd__or2_1
XFILLER_53_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09313_ _11507_/Q _09293_/X _09312_/X vssd1 vssd1 vccd1 vccd1 _11507_/D sky130_fd_sc_hd__a21o_1
XFILLER_146_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06525_ _11707_/Q _08560_/A _06522_/X _06524_/X vssd1 vssd1 vccd1 vccd1 _06525_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09244_ _09243_/B _07037_/B _09229_/Y _09243_/X vssd1 vssd1 vccd1 vccd1 _11474_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_139_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06456_ _10426_/Q _06541_/A2 _06504_/B1 _11008_/Q _06455_/X vssd1 vssd1 vccd1 vccd1
+ _06456_/X sky130_fd_sc_hd__o221a_1
XFILLER_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05407_ _10582_/Q _10581_/Q _05418_/S vssd1 vssd1 vccd1 vccd1 _05411_/A sky130_fd_sc_hd__mux2_1
X_09175_ _09226_/A _09175_/B vssd1 vssd1 vccd1 vccd1 _09175_/Y sky130_fd_sc_hd__nor2_2
X_06387_ _06387_/A _06387_/B _06387_/C vssd1 vssd1 vccd1 vccd1 _06387_/X sky130_fd_sc_hd__and3_2
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08126_ _08579_/A0 _10889_/Q _08140_/S vssd1 vssd1 vccd1 vccd1 _08127_/B sky130_fd_sc_hd__mux2_1
X_05338_ _11094_/Q _11093_/Q _05426_/S vssd1 vssd1 vccd1 vccd1 _05340_/C sky130_fd_sc_hd__mux2_1
X_08057_ _10854_/Q _08426_/B vssd1 vssd1 vccd1 vccd1 _08057_/X sky130_fd_sc_hd__or2_1
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05269_ _05269_/A _05269_/B _05269_/C _05269_/D vssd1 vssd1 vccd1 vccd1 _05270_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_135_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07008_ _07617_/A _07090_/A vssd1 vssd1 vccd1 vccd1 _07008_/X sky130_fd_sc_hd__or2_4
XFILLER_89_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput104 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 input104/X sky130_fd_sc_hd__buf_4
Xinput115 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 input115/X sky130_fd_sc_hd__buf_6
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08959_ _09538_/B _09539_/A _09668_/A vssd1 vssd1 vccd1 vccd1 _08959_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10921_ _11220_/CLK _10921_/D vssd1 vssd1 vccd1 vccd1 _10921_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10852_ _11641_/CLK _10852_/D vssd1 vssd1 vccd1 vccd1 _10852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _11472_/CLK _10783_/D vssd1 vssd1 vccd1 vccd1 _10783_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11404_ _11495_/CLK _11404_/D vssd1 vssd1 vccd1 vccd1 _11404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11335_ _11756_/CLK _11335_/D vssd1 vssd1 vccd1 vccd1 _11335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11266_ _11268_/CLK _11266_/D vssd1 vssd1 vccd1 vccd1 _11266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10217_ _11634_/CLK _10217_/D vssd1 vssd1 vccd1 vccd1 _10217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11197_ _11251_/CLK _11197_/D vssd1 vssd1 vccd1 vccd1 _11197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10148_ _11787_/Q _10154_/B vssd1 vssd1 vccd1 vccd1 _10148_/X sky130_fd_sc_hd__or2_1
XFILLER_132_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10079_ _10115_/A0 _11739_/Q _10082_/S vssd1 vssd1 vccd1 vccd1 _11739_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06310_ _06300_/X _06301_/X _06304_/X _06309_/X vssd1 vssd1 vccd1 vccd1 _06310_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_91_1368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07290_ _07936_/A _07290_/B vssd1 vssd1 vccd1 vccd1 _10413_/D sky130_fd_sc_hd__or2_1
X_06241_ _10751_/Q _07853_/A _07540_/A _10561_/Q vssd1 vssd1 vccd1 vccd1 _06241_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_50_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06172_ _11544_/Q _09359_/A _06168_/X _06171_/X vssd1 vssd1 vccd1 vccd1 _06178_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05123_ _05123_/A _05123_/B _05123_/C _05123_/D vssd1 vssd1 vccd1 vccd1 _05124_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09931_ _11663_/Q _09851_/Y _09908_/Y _06955_/X _09930_/Y vssd1 vssd1 vccd1 vccd1
+ _09931_/X sky130_fd_sc_hd__a221o_1
Xfanout805 _06166_/A2 vssd1 vssd1 vccd1 vccd1 _06351_/A2 sky130_fd_sc_hd__buf_6
Xfanout816 _06735_/B1 vssd1 vssd1 vccd1 vccd1 _09038_/A sky130_fd_sc_hd__buf_8
XFILLER_131_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout827 _06238_/A2 vssd1 vssd1 vccd1 vccd1 _07190_/A sky130_fd_sc_hd__buf_8
X_09862_ _11444_/Q _09881_/A2 _09881_/B1 _10703_/Q vssd1 vssd1 vccd1 vccd1 _09868_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout838 fanout846/X vssd1 vssd1 vccd1 vccd1 _06803_/A2 sky130_fd_sc_hd__buf_6
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout849 _05742_/Y vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__buf_12
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _08819_/A _08813_/B vssd1 vssd1 vccd1 vccd1 _11263_/D sky130_fd_sc_hd__or2_1
XFILLER_140_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _11650_/Q _09404_/Y _09792_/X _09681_/B vssd1 vssd1 vccd1 vccd1 _09793_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05956_ _11541_/Q _06219_/A2 _05952_/X _05955_/X vssd1 vssd1 vccd1 vccd1 _05962_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08744_ _08834_/A0 _11229_/Q _08748_/S vssd1 vssd1 vccd1 vccd1 _08745_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _09985_/A1 _11192_/Q _08695_/S vssd1 vssd1 vccd1 vccd1 _08676_/B sky130_fd_sc_hd__mux2_1
X_05887_ _11520_/Q _09326_/A _06363_/A2 _11480_/Q vssd1 vssd1 vccd1 vccd1 _05887_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07626_ _07316_/X _10598_/Q _07626_/S vssd1 vssd1 vccd1 vccd1 _10598_/D sky130_fd_sc_hd__mux2_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07557_ _09289_/A1 _10562_/Q _07557_/S vssd1 vssd1 vccd1 vccd1 _07558_/B sky130_fd_sc_hd__mux2_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06508_ _10849_/Q _06643_/A2 _06642_/A2 _10470_/Q _06507_/X vssd1 vssd1 vccd1 vccd1
+ _06508_/X sky130_fd_sc_hd__o221a_1
XFILLER_10_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07488_ _07093_/X _10524_/Q _07491_/S vssd1 vssd1 vccd1 vccd1 _10524_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06439_ _10689_/Q _09358_/A _09976_/A _10511_/Q _06651_/C1 vssd1 vssd1 vccd1 vccd1
+ _06439_/X sky130_fd_sc_hd__a221o_1
X_09227_ _09227_/A _09243_/C vssd1 vssd1 vccd1 vccd1 _09227_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09158_ _11423_/Q _09154_/X _09157_/X vssd1 vssd1 vccd1 vccd1 _11423_/D sky130_fd_sc_hd__a21o_1
XFILLER_148_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08109_ _08193_/A _08109_/B vssd1 vssd1 vccd1 vccd1 _10879_/D sky130_fd_sc_hd__or2_1
X_09089_ _11392_/Q _09099_/B vssd1 vssd1 vccd1 vccd1 _09089_/X sky130_fd_sc_hd__or2_1
XFILLER_107_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11120_ _11812_/CLK _11120_/D vssd1 vssd1 vccd1 vccd1 _11120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _11291_/CLK _11051_/D vssd1 vssd1 vccd1 vccd1 _11051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10002_ _10112_/A0 _11689_/Q _10008_/S vssd1 vssd1 vccd1 vccd1 _11689_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10904_ _11284_/CLK _10904_/D vssd1 vssd1 vccd1 vccd1 _10904_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ _11657_/CLK _10835_/D vssd1 vssd1 vccd1 vccd1 _10835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10766_ _11439_/CLK _10766_/D vssd1 vssd1 vccd1 vccd1 _10766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ _11573_/CLK _10697_/D vssd1 vssd1 vccd1 vccd1 _10697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _11411_/CLK _11318_/D vssd1 vssd1 vccd1 vccd1 _11318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11249_ _11572_/CLK _11249_/D vssd1 vssd1 vccd1 vccd1 _11249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05810_ _10935_/Q _06630_/A2 _06630_/B1 _11011_/Q vssd1 vssd1 vccd1 vccd1 _05810_/X
+ sky130_fd_sc_hd__o22a_1
X_06790_ _10413_/Q _06804_/B vssd1 vssd1 vccd1 vccd1 _06790_/X sky130_fd_sc_hd__or2_1
XFILLER_110_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05741_ _05751_/B _05749_/A _05745_/A vssd1 vssd1 vccd1 vccd1 _05741_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_76_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08460_ _08821_/A _08460_/B vssd1 vssd1 vccd1 vccd1 _11080_/D sky130_fd_sc_hd__and2_1
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05672_ _11197_/Q _05549_/Y _05603_/Y _11193_/Q vssd1 vssd1 vccd1 vccd1 _05679_/C
+ sky130_fd_sc_hd__a22o_1
X_07411_ _09214_/A _10482_/Q _07425_/S vssd1 vssd1 vccd1 vccd1 _07412_/B sky130_fd_sc_hd__mux2_1
XFILLER_63_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08391_ _09985_/A1 _08414_/S _08390_/X _08791_/C1 vssd1 vssd1 vccd1 vccd1 _11036_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07342_ _10438_/Q _07350_/S _07346_/B1 _07227_/B vssd1 vssd1 vccd1 vccd1 _10438_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_91_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07273_ _10405_/Q _09175_/B vssd1 vssd1 vccd1 vccd1 _07273_/X sky130_fd_sc_hd__or2_1
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _11357_/Q _08994_/X _09011_/X vssd1 vssd1 vccd1 vccd1 _11357_/D sky130_fd_sc_hd__a21o_1
X_06224_ _11763_/Q _10108_/A _08311_/A _10998_/Q vssd1 vssd1 vccd1 vccd1 _06224_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06155_ _11129_/Q _06635_/A2 _06514_/A2 _11261_/Q _06154_/X vssd1 vssd1 vccd1 vccd1
+ _06155_/X sky130_fd_sc_hd__o221a_1
XFILLER_105_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05106_ _11264_/Q _11263_/Q _05394_/S vssd1 vssd1 vccd1 vccd1 _05107_/D sky130_fd_sc_hd__mux2_1
X_06086_ _11543_/Q _06219_/A2 _06084_/X _06085_/X vssd1 vssd1 vccd1 vccd1 _06086_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout602 _08166_/A vssd1 vssd1 vccd1 vccd1 _06591_/A2 sky130_fd_sc_hd__clkbuf_8
X_09914_ _10484_/Q _09573_/B _09571_/D _10479_/Q _09913_/X vssd1 vssd1 vccd1 vccd1
+ _09917_/C sky130_fd_sc_hd__a221o_1
XFILLER_28_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout613 _06318_/A2 vssd1 vssd1 vccd1 vccd1 _06541_/A2 sky130_fd_sc_hd__buf_4
Xfanout624 _06735_/A2 vssd1 vssd1 vccd1 vccd1 _09060_/A sky130_fd_sc_hd__buf_8
XFILLER_28_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout635 _09833_/A vssd1 vssd1 vccd1 vccd1 _09529_/A sky130_fd_sc_hd__buf_4
XFILLER_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout646 _05619_/A1 vssd1 vssd1 vccd1 vccd1 _05631_/A2 sky130_fd_sc_hd__buf_6
Xfanout657 _11628_/Q vssd1 vssd1 vccd1 vccd1 _05629_/A2 sky130_fd_sc_hd__buf_6
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _11460_/Q _09879_/A2 _09886_/B1 _10786_/Q _09844_/X vssd1 vssd1 vccd1 vccd1
+ _09850_/B sky130_fd_sc_hd__a221o_1
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout668 _09430_/B vssd1 vssd1 vccd1 vccd1 _09680_/B sky130_fd_sc_hd__buf_8
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout679 _05413_/S vssd1 vssd1 vccd1 vccd1 _05430_/S sky130_fd_sc_hd__buf_12
XFILLER_86_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09776_ _09775_/B _09775_/C _11652_/Q vssd1 vssd1 vccd1 vccd1 _09776_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06988_ _10149_/A1 _06976_/X _06987_/X _06996_/C1 vssd1 vssd1 vccd1 vccd1 _10261_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _08821_/A _08727_/B vssd1 vssd1 vccd1 vccd1 _11220_/D sky130_fd_sc_hd__and2_1
XFILLER_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05939_ _11025_/Q _06629_/A2 _05935_/X _05938_/X vssd1 vssd1 vccd1 vccd1 _05939_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _07232_/B _08750_/B _08657_/X vssd1 vssd1 vccd1 vccd1 _11184_/D sky130_fd_sc_hd__a21o_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _10589_/Q _07597_/Y _07600_/Y _07316_/X vssd1 vssd1 vccd1 vccd1 _10589_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08589_ _08838_/A0 _11150_/Q _08589_/S vssd1 vssd1 vccd1 vccd1 _08590_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ _11766_/CLK _10620_/D vssd1 vssd1 vccd1 vccd1 _10620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10551_ _10785_/CLK _10551_/D vssd1 vssd1 vccd1 vccd1 _10551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10482_ _11661_/CLK _10482_/D vssd1 vssd1 vccd1 vccd1 _10482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11103_ _11411_/CLK _11103_/D vssd1 vssd1 vccd1 vccd1 _11103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11034_ _11393_/CLK _11034_/D vssd1 vssd1 vccd1 vccd1 _11034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _11867_/A vssd1 vssd1 vccd1 vccd1 _11867_/X sky130_fd_sc_hd__buf_2
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10818_ _11584_/CLK _10818_/D vssd1 vssd1 vccd1 vccd1 _10818_/Q sky130_fd_sc_hd__dfxtp_1
X_11798_ _11800_/CLK _11798_/D vssd1 vssd1 vccd1 vccd1 _11798_/Q sky130_fd_sc_hd__dfxtp_1
X_10749_ _11622_/CLK _10749_/D vssd1 vssd1 vccd1 vccd1 _10749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput205 _05480_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07960_ _07037_/X _10802_/Q _07961_/S vssd1 vssd1 vccd1 vccd1 _10802_/D sky130_fd_sc_hd__mux2_1
X_06911_ _09256_/A1 _06903_/X _06910_/X _06990_/C1 vssd1 vssd1 vccd1 vccd1 _10196_/D
+ sky130_fd_sc_hd__o211a_1
X_07891_ _10764_/Q _07901_/B vssd1 vssd1 vccd1 vccd1 _07891_/X sky130_fd_sc_hd__or2_1
X_09630_ _10729_/Q _09565_/A _09573_/D _10720_/Q _09621_/X vssd1 vssd1 vccd1 vccd1
+ _09633_/B sky130_fd_sc_hd__a221o_1
X_06842_ _11448_/Q _07777_/A _07254_/A _10415_/Q vssd1 vssd1 vccd1 vccd1 _06842_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06773_ _10528_/Q _06873_/A2 _06710_/B _10733_/Q _06772_/X vssd1 vssd1 vccd1 vccd1
+ _06773_/X sky130_fd_sc_hd__o221a_1
XFILLER_3_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09561_ _09600_/B _09561_/B vssd1 vssd1 vccd1 vccd1 _09823_/A sky130_fd_sc_hd__nor2_2
XFILLER_23_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08512_ _08783_/A _08512_/B vssd1 vssd1 vccd1 vccd1 _11105_/D sky130_fd_sc_hd__or2_1
XFILLER_36_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05724_ _10973_/Q _05591_/Y _05633_/Y _10956_/Q vssd1 vssd1 vccd1 vccd1 _05724_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09492_ _09528_/B _09492_/B _09489_/B vssd1 vssd1 vccd1 vccd1 _09492_/X sky130_fd_sc_hd__or3b_1
XFILLER_97_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08443_ _11064_/Q _08437_/Y _08438_/Y _07314_/X vssd1 vssd1 vccd1 vccd1 _11064_/D
+ sky130_fd_sc_hd__o22a_1
X_05655_ _05655_/A _05655_/B _05655_/C _05655_/D vssd1 vssd1 vccd1 vccd1 _05655_/X
+ sky130_fd_sc_hd__or4_2
X_08374_ _11029_/Q _08438_/B vssd1 vssd1 vccd1 vccd1 _08374_/X sky130_fd_sc_hd__or2_1
X_05586_ _05628_/A2 _10200_/Q _10197_/Q _05628_/B1 vssd1 vssd1 vccd1 vccd1 _05586_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07325_ _07599_/A _08164_/B vssd1 vssd1 vccd1 vccd1 _07325_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07256_ _07818_/A _07256_/B vssd1 vssd1 vccd1 vccd1 _10396_/D sky130_fd_sc_hd__or2_1
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06207_ _06633_/A _06162_/X _06167_/X _06619_/A1 _06157_/X vssd1 vssd1 vccd1 vccd1
+ _06207_/X sky130_fd_sc_hd__o311a_2
X_07187_ _09214_/B _07187_/B vssd1 vssd1 vccd1 vccd1 _07187_/X sky130_fd_sc_hd__or2_1
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06138_ _10789_/Q _06540_/A2 _06538_/B1 _10638_/Q vssd1 vssd1 vccd1 vccd1 _06138_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06069_ _11027_/Q _06538_/A2 _06065_/X _06068_/X vssd1 vssd1 vccd1 vccd1 _06075_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout410 _05368_/Y vssd1 vssd1 vccd1 vccd1 _09944_/B1 sky130_fd_sc_hd__buf_8
Xfanout421 _05313_/Y vssd1 vssd1 vccd1 vccd1 _09876_/B1 sky130_fd_sc_hd__buf_6
XFILLER_132_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout432 _05248_/Y vssd1 vssd1 vccd1 vccd1 _09566_/C sky130_fd_sc_hd__buf_8
XFILLER_63_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout443 _05190_/Y vssd1 vssd1 vccd1 vccd1 _09873_/A2 sky130_fd_sc_hd__buf_4
Xfanout454 _05124_/Y vssd1 vssd1 vccd1 vccd1 _09567_/A sky130_fd_sc_hd__buf_6
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout465 _08588_/C1 vssd1 vssd1 vccd1 vccd1 _08345_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout476 _10153_/C1 vssd1 vssd1 vccd1 vccd1 _10155_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09828_ _09497_/A _09824_/S _09825_/A vssd1 vssd1 vccd1 vccd1 _09828_/Y sky130_fd_sc_hd__o21ai_1
Xfanout487 _07866_/C1 vssd1 vssd1 vccd1 vccd1 _07884_/C1 sky130_fd_sc_hd__buf_4
XFILLER_74_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout498 fanout510/X vssd1 vssd1 vccd1 vccd1 _09168_/C1 sky130_fd_sc_hd__buf_4
XFILLER_100_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09759_ _09515_/C _09722_/Y _09758_/Y _06948_/X vssd1 vssd1 vccd1 vccd1 _09759_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _11722_/CLK _11721_/D vssd1 vssd1 vccd1 vccd1 _11721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11652_/CLK _11652_/D vssd1 vssd1 vccd1 vccd1 _11652_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10603_ _11777_/CLK _10603_/D vssd1 vssd1 vccd1 vccd1 _10603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11583_ _11584_/CLK _11583_/D vssd1 vssd1 vccd1 vccd1 _11583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10534_ _10805_/CLK _10534_/D vssd1 vssd1 vccd1 vccd1 _10534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10465_ _10981_/CLK _10465_/D vssd1 vssd1 vccd1 vccd1 _10465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10396_ _10765_/CLK _10396_/D vssd1 vssd1 vccd1 vccd1 _10396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11017_ _11023_/CLK _11017_/D vssd1 vssd1 vccd1 vccd1 _11017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_66_wb_clk_i clkbuf_leaf_69_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11801_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1090 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1090/HI io_oeb[20] sky130_fd_sc_hd__conb_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05440_ _10678_/Q _09572_/C _09572_/D _10661_/Q vssd1 vssd1 vccd1 vccd1 _05440_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05371_ _10823_/Q _10822_/Q _05429_/S vssd1 vssd1 vccd1 vccd1 _05373_/C sky130_fd_sc_hd__mux2_1
X_07110_ _07111_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _07110_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08090_ _07005_/A _08091_/C _08089_/X vssd1 vssd1 vccd1 vccd1 _10870_/D sky130_fd_sc_hd__a21o_1
XFILLER_88_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07041_ _10278_/Q _07040_/X _07044_/S vssd1 vssd1 vccd1 vccd1 _10278_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _11348_/Q _08972_/X _08991_/X vssd1 vssd1 vccd1 vccd1 _11348_/D sky130_fd_sc_hd__a21o_1
XFILLER_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07943_ _08438_/A _08085_/B vssd1 vssd1 vccd1 vccd1 _07943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07874_ _08883_/A1 _07970_/S _07873_/X _07894_/C1 vssd1 vssd1 vccd1 vccd1 _10755_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09613_ _10628_/Q _09572_/B _09572_/C _10394_/Q _09610_/X vssd1 vssd1 vccd1 vccd1
+ _09615_/C sky130_fd_sc_hd__a221o_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06825_ _06852_/A1 _10247_/Q _06853_/A3 _06824_/X _05819_/B vssd1 vssd1 vccd1 vccd1
+ _06825_/X sky130_fd_sc_hd__a32o_1
XFILLER_37_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _11624_/Q _09541_/Y _09543_/X _09833_/A vssd1 vssd1 vccd1 vccd1 _11624_/D
+ sky130_fd_sc_hd__o211a_1
X_06756_ _11620_/Q _06704_/B _06755_/X vssd1 vssd1 vccd1 vccd1 _10242_/D sky130_fd_sc_hd__a21o_1
XFILLER_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05707_ _11036_/Q _05567_/Y _05621_/Y _11045_/Q vssd1 vssd1 vccd1 vccd1 _05709_/C
+ sky130_fd_sc_hd__a22o_1
X_06687_ _10488_/Q _06872_/A2 _06710_/B _10799_/Q vssd1 vssd1 vccd1 vccd1 _06687_/X
+ sky130_fd_sc_hd__o22a_1
X_09475_ _09475_/A _09475_/B vssd1 vssd1 vccd1 vccd1 _09475_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08426_ _08438_/A _08426_/B vssd1 vssd1 vccd1 vccd1 _08426_/Y sky130_fd_sc_hd__nor2_2
X_05638_ _11326_/Q _05615_/Y _05621_/Y _11325_/Q _05637_/X vssd1 vssd1 vccd1 vccd1
+ _05643_/A sky130_fd_sc_hd__a221o_1
XFILLER_145_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05569_ _05618_/A1 _11415_/Q _11412_/Q _05606_/B2 vssd1 vssd1 vccd1 vccd1 _05569_/X
+ sky130_fd_sc_hd__a22o_1
X_08357_ _08839_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _11021_/D sky130_fd_sc_hd__or2_1
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07308_ _10419_/Q _07301_/Y _07306_/Y _07229_/X vssd1 vssd1 vccd1 vccd1 _10419_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08288_ _08745_/A _08467_/S vssd1 vssd1 vccd1 vccd1 _08298_/S sky130_fd_sc_hd__or2_4
XFILLER_125_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07239_ _07025_/A _07665_/S _07928_/A vssd1 vssd1 vccd1 vccd1 _07239_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10250_ _10769_/CLK _10250_/D vssd1 vssd1 vccd1 vccd1 _10250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10181_ _10181_/A0 _11802_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _11802_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout240 _09491_/X vssd1 vssd1 vccd1 vccd1 _09528_/B sky130_fd_sc_hd__buf_4
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout251 _08765_/X vssd1 vssd1 vccd1 vccd1 _08792_/S sky130_fd_sc_hd__buf_6
Xfanout262 _08472_/X vssd1 vssd1 vccd1 vccd1 _08497_/S sky130_fd_sc_hd__buf_4
Xfanout273 _08166_/X vssd1 vssd1 vccd1 vccd1 _08182_/S sky130_fd_sc_hd__buf_4
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout284 _07890_/A2 vssd1 vssd1 vccd1 vccd1 _07871_/S sky130_fd_sc_hd__buf_6
Xfanout295 _07778_/X vssd1 vssd1 vccd1 vccd1 _09200_/S sky130_fd_sc_hd__buf_8
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11706_/CLK _11704_/D vssd1 vssd1 vccd1 vccd1 _11704_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ _11652_/CLK _11635_/D vssd1 vssd1 vccd1 vccd1 _11635_/Q sky130_fd_sc_hd__dfxtp_1
X_11566_ _11758_/CLK _11566_/D vssd1 vssd1 vccd1 vccd1 _11566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10517_ _11474_/CLK _10517_/D vssd1 vssd1 vccd1 vccd1 _10517_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11497_ _11497_/CLK _11497_/D vssd1 vssd1 vccd1 vccd1 _11497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_113_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11474_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10448_ _11777_/CLK _10448_/D vssd1 vssd1 vccd1 vccd1 _10448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10379_ _10812_/CLK _10379_/D vssd1 vssd1 vccd1 vccd1 _10379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06610_ _10486_/Q _08649_/A _06608_/X _06609_/X vssd1 vssd1 vccd1 vccd1 _06610_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07590_ _07796_/A _07590_/B vssd1 vssd1 vccd1 vccd1 _10578_/D sky130_fd_sc_hd__or2_1
XFILLER_20_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06541_ _11236_/Q _06541_/A2 _06589_/A2 _11010_/Q _06540_/X vssd1 vssd1 vccd1 vccd1
+ _06541_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ _10149_/A1 _09266_/B _08761_/A vssd1 vssd1 vccd1 vccd1 _09260_/X sky130_fd_sc_hd__a21o_1
X_06472_ _10619_/Q _06642_/A2 _06471_/X _07083_/B vssd1 vssd1 vccd1 vccd1 _06472_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05423_ _05423_/A _05423_/B vssd1 vssd1 vccd1 vccd1 _05423_/Y sky130_fd_sc_hd__nor2_8
X_08211_ _10114_/A0 _10940_/Q _08219_/S vssd1 vssd1 vccd1 vccd1 _08212_/B sky130_fd_sc_hd__mux2_1
X_09191_ _09227_/A _09193_/B vssd1 vssd1 vccd1 vccd1 _09191_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05354_ _05354_/A _05354_/B _05354_/C _05354_/D vssd1 vssd1 vccd1 vccd1 _05357_/A
+ sky130_fd_sc_hd__or4_4
X_08142_ _08834_/A0 _10897_/Q _08146_/S vssd1 vssd1 vccd1 vccd1 _08143_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08073_ _10862_/Q _08085_/B vssd1 vssd1 vccd1 vccd1 _08073_/X sky130_fd_sc_hd__or2_1
XFILLER_146_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05285_ _10890_/Q _10889_/Q _05429_/S vssd1 vssd1 vccd1 vccd1 _05290_/B sky130_fd_sc_hd__mux2_1
X_07024_ _10134_/A0 _07000_/B _07000_/Y _10272_/Q _07309_/A vssd1 vssd1 vccd1 vccd1
+ _10272_/D sky130_fd_sc_hd__a221o_1
XFILLER_31_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08975_ _09275_/A1 _08989_/B _09290_/B1 vssd1 vssd1 vccd1 vccd1 _08975_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07926_ _07926_/A _07926_/B vssd1 vssd1 vccd1 vccd1 _10780_/D sky130_fd_sc_hd__or2_1
XFILLER_64_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07857_ _10747_/Q _07883_/B vssd1 vssd1 vccd1 vccd1 _07857_/X sky130_fd_sc_hd__or2_1
XFILLER_72_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06808_ _11459_/Q _06862_/A2 _06807_/X _06808_/C1 vssd1 vssd1 vccd1 vccd1 _06808_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07788_ _08536_/A _07788_/B vssd1 vssd1 vccd1 vccd1 _10701_/D sky130_fd_sc_hd__or2_1
XFILLER_25_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09527_ _09502_/A _09489_/C _09500_/C _11619_/Q vssd1 vssd1 vccd1 vccd1 _09529_/B
+ sky130_fd_sc_hd__a31o_1
X_06739_ _11304_/Q _06739_/A2 _06735_/X _06738_/X vssd1 vssd1 vccd1 vccd1 _06739_/X
+ sky130_fd_sc_hd__o211a_2
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _05426_/S _09475_/A _09457_/Y _09407_/A vssd1 vssd1 vccd1 vccd1 _11597_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08409_ _08793_/A _08409_/B vssd1 vssd1 vccd1 vccd1 _11045_/D sky130_fd_sc_hd__or2_1
XFILLER_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09389_ _10105_/A1 _11556_/Q _09390_/S vssd1 vssd1 vccd1 vccd1 _11556_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11420_ _11792_/CLK _11420_/D vssd1 vssd1 vccd1 vccd1 _11420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11351_ _11811_/CLK _11351_/D vssd1 vssd1 vccd1 vccd1 _11351_/Q sky130_fd_sc_hd__dfxtp_1
X_10302_ _11776_/CLK _10302_/D vssd1 vssd1 vccd1 vccd1 _10302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ _11284_/CLK _11282_/D vssd1 vssd1 vccd1 vccd1 _11282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10233_ _11702_/CLK _10233_/D vssd1 vssd1 vccd1 vccd1 _10233_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10164_ _11794_/Q _10176_/B vssd1 vssd1 vccd1 vccd1 _10164_/X sky130_fd_sc_hd__or2_1
Xfanout1002 input81/X vssd1 vssd1 vccd1 vccd1 _11868_/A sky130_fd_sc_hd__buf_6
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1013 input117/X vssd1 vssd1 vccd1 vccd1 _09129_/A1 sky130_fd_sc_hd__buf_12
Xfanout1024 _07018_/A vssd1 vssd1 vccd1 vccd1 _10080_/A0 sky130_fd_sc_hd__buf_4
Xfanout1035 _10172_/A1 vssd1 vssd1 vccd1 vccd1 _09124_/A1 sky130_fd_sc_hd__buf_4
XFILLER_86_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1046 _09396_/A0 vssd1 vssd1 vccd1 vccd1 _10113_/A0 sky130_fd_sc_hd__buf_4
X_10095_ _10184_/A0 _10087_/X _10094_/X _10155_/C1 vssd1 vssd1 vccd1 vccd1 _11749_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout1057 _07010_/A vssd1 vssd1 vccd1 vccd1 _10184_/A0 sky130_fd_sc_hd__buf_6
XFILLER_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1068 _10165_/A1 vssd1 vssd1 vccd1 vccd1 _09276_/A1 sky130_fd_sc_hd__buf_6
Xfanout1079 input100/X vssd1 vssd1 vccd1 vccd1 _07932_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10997_ _11763_/CLK _10997_/D vssd1 vssd1 vccd1 vccd1 _10997_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ _11622_/CLK _11618_/D vssd1 vssd1 vccd1 vccd1 _11618_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11549_ _11758_/CLK _11549_/D vssd1 vssd1 vccd1 vccd1 _11549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08760_ _08760_/A0 _11237_/Q _08760_/S vssd1 vssd1 vccd1 vccd1 _08761_/B sky130_fd_sc_hd__mux2_1
X_05972_ _10206_/Q _06351_/A2 _05968_/X _05971_/X vssd1 vssd1 vccd1 vccd1 _05972_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_wb_clk_i clkbuf_leaf_85_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11573_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07711_ _07785_/A0 _07755_/A2 _07710_/X _07866_/C1 vssd1 vssd1 vccd1 vccd1 _10656_/D
+ sky130_fd_sc_hd__o211a_1
X_08691_ _08789_/A1 _11200_/Q _08695_/S vssd1 vssd1 vccd1 vccd1 _08692_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11140_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07642_ _08901_/A1 _10609_/Q _07642_/S vssd1 vssd1 vccd1 vccd1 _10609_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07573_ _07025_/A _10570_/Q _07593_/S vssd1 vssd1 vccd1 vccd1 _07574_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09312_ _10178_/A1 _09310_/B _10178_/B1 vssd1 vssd1 vccd1 vccd1 _09312_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06524_ _10690_/Q _09358_/A _09976_/A _10513_/Q _07151_/A vssd1 vssd1 vccd1 vccd1
+ _06524_/X sky130_fd_sc_hd__a221o_1
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09243_ _11474_/Q _09243_/B _09243_/C vssd1 vssd1 vccd1 vccd1 _09243_/X sky130_fd_sc_hd__and3_1
XFILLER_146_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06455_ _10866_/Q _06455_/A2 _06455_/B1 _10432_/Q vssd1 vssd1 vccd1 vccd1 _06455_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05406_ _05406_/A _05406_/B _05406_/C _05406_/D vssd1 vssd1 vccd1 vccd1 _05412_/A
+ sky130_fd_sc_hd__or4_2
X_09174_ _11431_/Q _09154_/X _09173_/X vssd1 vssd1 vccd1 vccd1 _11431_/D sky130_fd_sc_hd__a21o_1
X_06386_ _10424_/Q _06541_/A2 _06504_/B1 _11006_/Q _06385_/X vssd1 vssd1 vccd1 vccd1
+ _06387_/C sky130_fd_sc_hd__o221a_1
XFILLER_147_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08125_ _09999_/A0 _08140_/S _08124_/X _08841_/C1 vssd1 vssd1 vccd1 vccd1 _10888_/D
+ sky130_fd_sc_hd__o211a_1
X_05337_ _11100_/Q _11099_/Q _05349_/S vssd1 vssd1 vccd1 vccd1 _05340_/B sky130_fd_sc_hd__mux2_1
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05268_ _10444_/Q _10739_/Q _05385_/S vssd1 vssd1 vccd1 vccd1 _05269_/D sky130_fd_sc_hd__mux2_1
X_08056_ _08835_/A _08056_/B vssd1 vssd1 vccd1 vccd1 _10853_/D sky130_fd_sc_hd__or2_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07007_ _07007_/A _10028_/A vssd1 vssd1 vccd1 vccd1 _07090_/A sky130_fd_sc_hd__and2_4
XFILLER_66_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05199_ _09539_/A _11026_/Q _05191_/X _05194_/X _05195_/X vssd1 vssd1 vccd1 vccd1
+ _05199_/X sky130_fd_sc_hd__a2111o_1
XFILLER_153_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput105 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 _07143_/A sky130_fd_sc_hd__buf_6
XFILLER_153_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput116 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 input116/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08958_ _08958_/A _09832_/S vssd1 vssd1 vccd1 vccd1 _08965_/A sky130_fd_sc_hd__nor2_2
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07909_ _10021_/A0 _10772_/Q _09206_/B vssd1 vssd1 vccd1 vccd1 _07910_/B sky130_fd_sc_hd__mux2_1
XFILLER_57_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08889_ _09216_/A0 _08884_/S _08888_/X _08943_/C1 vssd1 vssd1 vccd1 vccd1 _11301_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10920_ _11770_/CLK _10920_/D vssd1 vssd1 vccd1 vccd1 _10920_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ _11641_/CLK _10851_/D vssd1 vssd1 vccd1 vccd1 _10851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10782_/CLK _10782_/D vssd1 vssd1 vccd1 vccd1 _10782_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11403_ _11411_/CLK _11403_/D vssd1 vssd1 vccd1 vccd1 _11403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11334_ _11657_/CLK _11334_/D vssd1 vssd1 vccd1 vccd1 _11334_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11265_ _11779_/CLK _11265_/D vssd1 vssd1 vccd1 vccd1 _11265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10216_ _10981_/CLK _10216_/D vssd1 vssd1 vccd1 vccd1 _10216_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11196_ _11329_/CLK _11196_/D vssd1 vssd1 vccd1 vccd1 _11196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _11786_/Q _10137_/X _10146_/X vssd1 vssd1 vccd1 vccd1 _11786_/D sky130_fd_sc_hd__a21o_1
XFILLER_43_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10078_ _10114_/A0 _11738_/Q _10082_/S vssd1 vssd1 vccd1 vccd1 _11738_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06240_ _11455_/Q _07904_/A vssd1 vssd1 vccd1 vccd1 _06240_/X sky130_fd_sc_hd__or2_1
XFILLER_54_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06171_ _11682_/Q _09977_/A _06169_/X _06170_/X vssd1 vssd1 vccd1 vccd1 _06171_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05122_ _10305_/Q _10304_/Q _05300_/S vssd1 vssd1 vccd1 vccd1 _05123_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09930_ _11663_/Q _09938_/B vssd1 vssd1 vccd1 vccd1 _09930_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout806 _06870_/B1 vssd1 vssd1 vccd1 vccd1 _06858_/B1 sky130_fd_sc_hd__buf_6
XFILLER_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _09861_/A _09861_/B _09861_/C _09861_/D vssd1 vssd1 vccd1 vccd1 _09869_/B
+ sky130_fd_sc_hd__or4_1
Xfanout817 _06735_/B1 vssd1 vssd1 vccd1 vccd1 _06221_/A2 sky130_fd_sc_hd__buf_4
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout828 fanout846/X vssd1 vssd1 vccd1 vccd1 _06238_/A2 sky130_fd_sc_hd__buf_6
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout839 _06861_/B vssd1 vssd1 vccd1 vccd1 _07854_/A sky130_fd_sc_hd__buf_6
X_08812_ _11263_/Q _10128_/A0 _08820_/S vssd1 vssd1 vccd1 vccd1 _08813_/B sky130_fd_sc_hd__mux2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _11651_/Q _09771_/Y _09791_/X _09554_/B _09406_/B vssd1 vssd1 vccd1 vccd1
+ _09792_/X sky130_fd_sc_hd__o221a_1
XFILLER_86_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08743_ _08745_/A _08743_/B vssd1 vssd1 vccd1 vccd1 _11228_/D sky130_fd_sc_hd__or2_1
X_05955_ _11679_/Q _08594_/A _05953_/X _05954_/X vssd1 vssd1 vccd1 vccd1 _05955_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08674_ _09276_/A1 _08695_/S _08673_/X _09168_/C1 vssd1 vssd1 vccd1 vccd1 _11191_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05886_ _06450_/A _10224_/Q vssd1 vssd1 vccd1 vccd1 _05886_/X sky130_fd_sc_hd__and2_1
XFILLER_148_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07625_ _07098_/X _10597_/Q _07628_/S vssd1 vssd1 vccd1 vccd1 _10597_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07556_ _08684_/A _07556_/B vssd1 vssd1 vccd1 vccd1 _10561_/D sky130_fd_sc_hd__or2_1
XFILLER_107_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06507_ _11229_/Q _08650_/A _06640_/B1 _11141_/Q vssd1 vssd1 vccd1 vccd1 _06507_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07487_ _07090_/X _10523_/Q _07490_/S vssd1 vssd1 vccd1 vccd1 _10523_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09226_ _09226_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09226_/Y sky130_fd_sc_hd__nor2_4
XFILLER_139_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06438_ _10288_/Q _09325_/A _09248_/A _10319_/Q vssd1 vssd1 vccd1 vccd1 _06438_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09157_ _10162_/A1 _09171_/B _09173_/B1 vssd1 vssd1 vccd1 vccd1 _09157_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06369_ _10344_/Q _07152_/A _06368_/X _06808_/C1 vssd1 vssd1 vccd1 vccd1 _06369_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08108_ _10879_/Q _07015_/A _08120_/S vssd1 vssd1 vccd1 vccd1 _08109_/B sky130_fd_sc_hd__mux2_1
X_09088_ _11391_/Q _09082_/X _09087_/X vssd1 vssd1 vccd1 vccd1 _11391_/D sky130_fd_sc_hd__a21o_1
X_08039_ _10844_/Q _07015_/A _08051_/S vssd1 vssd1 vccd1 vccd1 _08040_/B sky130_fd_sc_hd__mux2_1
XFILLER_150_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11050_ _11812_/CLK _11050_/D vssd1 vssd1 vccd1 vccd1 _11050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10001_ _10111_/A0 _11688_/Q _10008_/S vssd1 vssd1 vccd1 vccd1 _11688_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903_ _11527_/CLK _10903_/D vssd1 vssd1 vccd1 vccd1 _10903_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10834_ _11243_/CLK _10834_/D vssd1 vssd1 vccd1 vccd1 _10834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10765_ _10765_/CLK _10765_/D vssd1 vssd1 vccd1 vccd1 _10765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10696_ _11711_/CLK _10696_/D vssd1 vssd1 vccd1 vccd1 _10696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11317_ _11330_/CLK _11317_/D vssd1 vssd1 vccd1 vccd1 _11317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11248_ _11319_/CLK _11248_/D vssd1 vssd1 vccd1 vccd1 _11248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11179_ _11268_/CLK _11179_/D vssd1 vssd1 vccd1 vccd1 _11179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05740_ _05751_/B _05749_/A _05745_/A vssd1 vssd1 vccd1 vccd1 _05740_/X sky130_fd_sc_hd__and3b_2
XFILLER_36_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05671_ _11206_/Q _05543_/Y _05615_/Y _11202_/Q vssd1 vssd1 vccd1 vccd1 _05679_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07410_ _07476_/A _07410_/B vssd1 vssd1 vccd1 vccd1 _10481_/D sky130_fd_sc_hd__or2_1
XFILLER_56_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08390_ _11036_/Q _08422_/B vssd1 vssd1 vccd1 vccd1 _08390_/X sky130_fd_sc_hd__or2_1
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07341_ _10437_/Q _07350_/S _07846_/S _07090_/A vssd1 vssd1 vccd1 vccd1 _10437_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_1343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07272_ _07928_/A _07272_/B vssd1 vssd1 vccd1 vccd1 _10404_/D sky130_fd_sc_hd__or2_1
XFILLER_143_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09011_ _10105_/A1 _09013_/B _08664_/A vssd1 vssd1 vccd1 vccd1 _09011_/X sky130_fd_sc_hd__a21o_1
X_06223_ _06218_/X _06219_/X _06222_/X _06217_/X vssd1 vssd1 vccd1 vccd1 _06223_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06154_ _10441_/Q _06513_/A2 _06126_/B _11213_/Q vssd1 vssd1 vccd1 vccd1 _06154_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_145_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05105_ _11260_/Q _11259_/Q _05393_/S vssd1 vssd1 vccd1 vccd1 _05107_/C sky130_fd_sc_hd__mux2_1
X_06085_ _11797_/Q _10159_/A _09293_/A _11503_/Q vssd1 vssd1 vccd1 vccd1 _06085_/X
+ sky130_fd_sc_hd__o22a_1
X_09913_ _10491_/Q _09573_/C _09950_/B1 _10483_/Q vssd1 vssd1 vccd1 vccd1 _09913_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout603 _06430_/A2 vssd1 vssd1 vccd1 vccd1 _08166_/A sky130_fd_sc_hd__buf_4
XFILLER_132_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout614 _07300_/A vssd1 vssd1 vccd1 vccd1 _06318_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout625 _06696_/A2 vssd1 vssd1 vccd1 vccd1 _06735_/A2 sky130_fd_sc_hd__buf_6
XFILLER_28_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout636 _09447_/B vssd1 vssd1 vccd1 vccd1 _09833_/A sky130_fd_sc_hd__buf_4
XFILLER_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout647 _05075_/Y vssd1 vssd1 vccd1 vccd1 _05619_/A1 sky130_fd_sc_hd__buf_8
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _10776_/Q _09884_/A2 _09565_/C _10778_/Q _09843_/X vssd1 vssd1 vccd1 vccd1
+ _09844_/X sky130_fd_sc_hd__a221o_1
XFILLER_59_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout658 _11628_/Q vssd1 vssd1 vccd1 vccd1 _09552_/A1 sky130_fd_sc_hd__buf_8
XFILLER_154_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout669 _11601_/Q vssd1 vssd1 vccd1 vccd1 _09430_/B sky130_fd_sc_hd__buf_12
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09775_ _11652_/Q _09775_/B _09775_/C vssd1 vssd1 vccd1 vccd1 _09775_/X sky130_fd_sc_hd__or3_1
X_06987_ _10261_/Q _06995_/B vssd1 vssd1 vccd1 vccd1 _06987_/X sky130_fd_sc_hd__or2_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ _11220_/Q _10135_/A0 _08726_/S vssd1 vssd1 vccd1 vccd1 _08727_/B sky130_fd_sc_hd__mux2_1
X_05938_ _10635_/Q _06453_/B1 _05937_/X _06265_/C1 vssd1 vssd1 vccd1 vccd1 _05938_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08657_ _11184_/Q _08437_/A _08742_/S _08303_/A vssd1 vssd1 vccd1 vccd1 _08657_/X
+ sky130_fd_sc_hd__a31o_1
X_05869_ _11124_/Q _06635_/A2 _05868_/X _06550_/C1 vssd1 vssd1 vccd1 vccd1 _05869_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _10588_/Q _07598_/Y _07599_/Y _07314_/X vssd1 vssd1 vccd1 vccd1 _10588_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08588_ _07107_/A _08589_/S _08587_/X _08588_/C1 vssd1 vssd1 vccd1 vccd1 _11149_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07539_ _07539_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07539_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10550_ _10773_/CLK _10550_/D vssd1 vssd1 vccd1 vccd1 _10550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09209_ _09229_/A _09221_/C vssd1 vssd1 vccd1 vccd1 _09209_/Y sky130_fd_sc_hd__nand2_4
XFILLER_10_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10481_ _11702_/CLK _10481_/D vssd1 vssd1 vccd1 vccd1 _10481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11102_ _11186_/CLK _11102_/D vssd1 vssd1 vccd1 vccd1 _11102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11033_ _11325_/CLK _11033_/D vssd1 vssd1 vccd1 vccd1 _11033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_138_wb_clk_i clkbuf_4_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11780_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ input79/X vssd1 vssd1 vccd1 vccd1 _11866_/X sky130_fd_sc_hd__buf_2
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10817_ _11310_/CLK _10817_/D vssd1 vssd1 vccd1 vccd1 _10817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11797_ _11801_/CLK _11797_/D vssd1 vssd1 vccd1 vccd1 _11797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10748_ _11442_/CLK _10748_/D vssd1 vssd1 vccd1 vccd1 _10748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10679_ _11458_/CLK _10679_/D vssd1 vssd1 vccd1 vccd1 _10679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput206 _05481_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_4
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06910_ _10196_/Q _06922_/B vssd1 vssd1 vccd1 vccd1 _06910_/X sky130_fd_sc_hd__or2_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07890_ input101/X _07890_/A2 _07889_/X _09201_/A1 vssd1 vssd1 vccd1 vccd1 _10763_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06841_ _10503_/Q _07440_/A vssd1 vssd1 vccd1 vccd1 _06841_/X sky130_fd_sc_hd__or2_1
XFILLER_96_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09560_ _11660_/Q _11645_/Q vssd1 vssd1 vccd1 vccd1 _09561_/B sky130_fd_sc_hd__nor2_2
X_06772_ _10393_/Q _06860_/A2 _06685_/B _11717_/Q vssd1 vssd1 vccd1 vccd1 _06772_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08511_ _09276_/A1 _11105_/Q _08537_/S vssd1 vssd1 vccd1 vccd1 _08512_/B sky130_fd_sc_hd__mux2_1
XFILLER_82_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05723_ _10958_/Q _05567_/Y _05621_/Y _10967_/Q vssd1 vssd1 vccd1 vccd1 _05727_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09491_ _09553_/A _09959_/B _09491_/C vssd1 vssd1 vccd1 vccd1 _09491_/X sky130_fd_sc_hd__or3_4
XFILLER_36_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08442_ _11063_/Q _08436_/Y _08439_/Y _09232_/B2 vssd1 vssd1 vccd1 vccd1 _11063_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05654_ _11301_/Q _05579_/Y _05597_/Y _11292_/Q _05645_/X vssd1 vssd1 vccd1 vccd1
+ _05655_/D sky130_fd_sc_hd__a221o_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08373_ _08757_/A _08373_/B vssd1 vssd1 vccd1 vccd1 _11028_/D sky130_fd_sc_hd__or2_1
X_05585_ _05585_/A _05585_/B vssd1 vssd1 vccd1 vccd1 _05585_/Y sky130_fd_sc_hd__nor2_8
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07324_ _07333_/A _07324_/B vssd1 vssd1 vccd1 vccd1 _07324_/X sky130_fd_sc_hd__or2_4
XFILLER_108_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07255_ _07303_/A _10396_/Q _09184_/S vssd1 vssd1 vccd1 vccd1 _07256_/B sky130_fd_sc_hd__mux2_1
X_06206_ _07151_/B _06200_/X _06205_/X _06189_/X vssd1 vssd1 vccd1 vccd1 _06206_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07186_ _07019_/X _10354_/Q _07186_/S vssd1 vssd1 vccd1 vccd1 _10354_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06137_ _10593_/Q _06539_/B1 _06455_/B1 _10903_/Q vssd1 vssd1 vccd1 vccd1 _06137_/X
+ sky130_fd_sc_hd__o22a_1
X_06068_ _10637_/Q _06538_/B1 _06067_/X _06265_/C1 vssd1 vssd1 vccd1 vccd1 _06068_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout400 _05423_/Y vssd1 vssd1 vccd1 vccd1 _09573_/D sky130_fd_sc_hd__buf_8
Xfanout411 _05368_/Y vssd1 vssd1 vccd1 vccd1 _09567_/D sky130_fd_sc_hd__buf_4
Xfanout422 _05302_/Y vssd1 vssd1 vccd1 vccd1 _09566_/D sky130_fd_sc_hd__buf_6
XFILLER_132_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout433 _05248_/Y vssd1 vssd1 vccd1 vccd1 _09886_/A2 sky130_fd_sc_hd__buf_4
XFILLER_99_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout444 _05179_/Y vssd1 vssd1 vccd1 vccd1 _09565_/A sky130_fd_sc_hd__buf_8
Xfanout455 _05124_/Y vssd1 vssd1 vccd1 vccd1 _09879_/A2 sky130_fd_sc_hd__buf_4
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout466 _08588_/C1 vssd1 vssd1 vccd1 vccd1 _08831_/C1 sky130_fd_sc_hd__buf_6
XFILLER_87_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09827_ _09827_/A _09827_/B vssd1 vssd1 vccd1 vccd1 _09827_/Y sky130_fd_sc_hd__xnor2_2
Xfanout477 _07018_/B vssd1 vssd1 vccd1 vccd1 _10153_/C1 sky130_fd_sc_hd__buf_4
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout488 _07882_/C1 vssd1 vssd1 vccd1 vccd1 _07866_/C1 sky130_fd_sc_hd__buf_4
XFILLER_74_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout499 _09048_/C1 vssd1 vssd1 vccd1 vccd1 _08937_/C1 sky130_fd_sc_hd__buf_4
XFILLER_41_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09758_ _09908_/A _09758_/B vssd1 vssd1 vccd1 vccd1 _09758_/Y sky130_fd_sc_hd__nor2_2
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08709_ _11209_/Q _07007_/A _08726_/S vssd1 vssd1 vccd1 vccd1 _08710_/B sky130_fd_sc_hd__mux2_1
XFILLER_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _11641_/Q _09692_/B vssd1 vssd1 vccd1 vccd1 _09689_/X sky130_fd_sc_hd__or2_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11720_/CLK _11720_/D vssd1 vssd1 vccd1 vccd1 _11720_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11651_/CLK _11651_/D vssd1 vssd1 vccd1 vccd1 _11651_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10602_ _11777_/CLK _10602_/D vssd1 vssd1 vccd1 vccd1 _10602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11582_ _11584_/CLK _11582_/D vssd1 vssd1 vccd1 vccd1 _11582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10533_ _10805_/CLK _10533_/D vssd1 vssd1 vccd1 vccd1 _10533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10464_ _10981_/CLK _10464_/D vssd1 vssd1 vccd1 vccd1 _10464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10395_ _11720_/CLK _10395_/D vssd1 vssd1 vccd1 vccd1 _10395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11016_ _11312_/CLK _11016_/D vssd1 vssd1 vccd1 vccd1 _11016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_tms1x00_1080 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1080/HI io_oeb[10] sky130_fd_sc_hd__conb_1
XFILLER_60_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1091 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1091/HI io_oeb[21] sky130_fd_sc_hd__conb_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05370_ _10872_/Q _10871_/Q _05426_/S vssd1 vssd1 vccd1 vccd1 _05373_/B sky130_fd_sc_hd__mux2_1
XFILLER_144_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11765_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07040_ _07451_/A _07040_/B vssd1 vssd1 vccd1 vccd1 _07040_/X sky130_fd_sc_hd__or2_4
XFILLER_146_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08991_ _09101_/A1 _08989_/B _09290_/B1 vssd1 vssd1 vccd1 vccd1 _08991_/X sky130_fd_sc_hd__a21o_1
XFILLER_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07942_ _08323_/A _08083_/S vssd1 vssd1 vccd1 vccd1 _07942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07873_ _10755_/Q _07893_/B vssd1 vssd1 vccd1 vccd1 _07873_/X sky130_fd_sc_hd__or2_1
XFILLER_96_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09612_ _10388_/Q _09565_/A _09573_/D _10383_/Q _09605_/X vssd1 vssd1 vccd1 vccd1
+ _09615_/B sky130_fd_sc_hd__a221o_1
X_06824_ _06852_/A1 _10247_/Q _06852_/A3 _06743_/X _06823_/X vssd1 vssd1 vccd1 vccd1
+ _06824_/X sky130_fd_sc_hd__a32o_1
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09543_ _11662_/Q _09538_/X _09542_/X vssd1 vssd1 vccd1 vccd1 _09543_/X sky130_fd_sc_hd__a21o_1
X_06755_ _06852_/A1 _10242_/Q _06853_/A3 _06754_/X _05819_/B vssd1 vssd1 vccd1 vccd1
+ _06755_/X sky130_fd_sc_hd__a32o_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05706_ _11041_/Q _05549_/Y _05603_/Y _11037_/Q vssd1 vssd1 vccd1 vccd1 _05709_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09474_ input39/X _09442_/X _09473_/X vssd1 vssd1 vccd1 vccd1 _09475_/B sky130_fd_sc_hd__o21ai_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06686_ _10692_/Q _07203_/A _06860_/A2 _10389_/Q _06685_/X vssd1 vssd1 vccd1 vccd1
+ _06686_/X sky130_fd_sc_hd__o221a_1
XFILLER_52_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08425_ _08437_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08425_/Y sky130_fd_sc_hd__nand2_2
XFILLER_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05637_ _11330_/Q _05543_/Y _05603_/Y _11317_/Q vssd1 vssd1 vccd1 vccd1 _05637_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08356_ _08834_/A0 _11021_/Q _08360_/S vssd1 vssd1 vccd1 vccd1 _08357_/B sky130_fd_sc_hd__mux2_1
X_05568_ _09552_/A1 _11420_/Q _11414_/Q _05078_/A vssd1 vssd1 vccd1 vccd1 _05568_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_138_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07307_ _10418_/Q _07301_/Y _07306_/Y _08326_/B2 vssd1 vssd1 vccd1 vccd1 _10418_/D
+ sky130_fd_sc_hd__a22o_1
X_08287_ _08745_/A _08467_/S vssd1 vssd1 vccd1 vccd1 _08287_/Y sky130_fd_sc_hd__nor2_1
X_05499_ _10244_/Q input56/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05499_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07238_ _10387_/Q _07246_/S _07237_/X _07012_/Y vssd1 vssd1 vccd1 vccd1 _10387_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07169_ _07796_/A _07169_/B vssd1 vssd1 vccd1 vccd1 _10345_/D sky130_fd_sc_hd__or2_1
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10180_ _10180_/A _10180_/B _10180_/C vssd1 vssd1 vccd1 vccd1 _10190_/S sky130_fd_sc_hd__or3_4
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout230 _07112_/Y vssd1 vssd1 vccd1 vccd1 _07188_/S sky130_fd_sc_hd__buf_8
Xfanout241 _09491_/X vssd1 vssd1 vccd1 vccd1 _09502_/B sky130_fd_sc_hd__buf_2
XFILLER_87_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout252 _08765_/X vssd1 vssd1 vccd1 vccd1 _08802_/S sky130_fd_sc_hd__buf_6
XFILLER_115_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout263 _08472_/X vssd1 vssd1 vccd1 vccd1 _08501_/S sky130_fd_sc_hd__buf_2
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout274 _08146_/S vssd1 vssd1 vccd1 vccd1 _08140_/S sky130_fd_sc_hd__buf_4
Xfanout285 _07890_/A2 vssd1 vssd1 vccd1 vccd1 _07970_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout296 _07645_/B vssd1 vssd1 vccd1 vccd1 _08197_/S sky130_fd_sc_hd__buf_6
XFILLER_47_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11703_/CLK _11703_/D vssd1 vssd1 vccd1 vccd1 _11703_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11634_/CLK _11634_/D vssd1 vssd1 vccd1 vccd1 _11634_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11565_ _11763_/CLK _11565_/D vssd1 vssd1 vccd1 vccd1 _11565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10516_ _10725_/CLK _10516_/D vssd1 vssd1 vccd1 vccd1 _10516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11496_ _11497_/CLK _11496_/D vssd1 vssd1 vccd1 vccd1 _11496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10447_ _11768_/CLK _10447_/D vssd1 vssd1 vccd1 vccd1 _10447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10378_ _11745_/CLK _10378_/D vssd1 vssd1 vccd1 vccd1 _10378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06540_ _10794_/Q _06540_/A2 _06540_/B1 _10434_/Q vssd1 vssd1 vccd1 vccd1 _06540_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06471_ _10461_/Q _06643_/A2 _08469_/B _10984_/Q _06470_/X vssd1 vssd1 vccd1 vccd1
+ _06471_/X sky130_fd_sc_hd__o221a_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_190 _07059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ _09396_/A0 _08219_/S _08209_/X _08351_/C1 vssd1 vssd1 vccd1 vccd1 _10939_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05422_ _05422_/A _05422_/B _05422_/C _05422_/D vssd1 vssd1 vccd1 vccd1 _05423_/B
+ sky130_fd_sc_hd__or4_4
X_09190_ _09226_/A _09192_/B vssd1 vssd1 vccd1 vccd1 _09190_/Y sky130_fd_sc_hd__nor2_4
XFILLER_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08141_ _08835_/A _08141_/B vssd1 vssd1 vccd1 vccd1 _10896_/D sky130_fd_sc_hd__or2_1
X_05353_ _11306_/Q _11305_/Q _05396_/S vssd1 vssd1 vccd1 vccd1 _05354_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08072_ _10088_/A1 _08083_/S _08071_/X _08662_/C1 vssd1 vssd1 vccd1 vccd1 _10861_/D
+ sky130_fd_sc_hd__o211a_1
X_05284_ _10898_/Q _10897_/Q _09680_/C vssd1 vssd1 vccd1 vccd1 _05290_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07023_ _10271_/Q _09232_/B2 _07038_/S vssd1 vssd1 vccd1 vccd1 _10271_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08974_ _09111_/A1 _08972_/X _08973_/X _09279_/C1 vssd1 vssd1 vccd1 vccd1 _11339_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07925_ _07028_/A _10780_/Q _09218_/S vssd1 vssd1 vccd1 vccd1 _07926_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07856_ _07303_/A _07970_/S _07855_/X _07894_/C1 vssd1 vssd1 vccd1 vccd1 _10746_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06807_ _10716_/Q _06807_/A2 _06861_/B _10765_/Q _06806_/X vssd1 vssd1 vccd1 vccd1
+ _06807_/X sky130_fd_sc_hd__o221a_2
XFILLER_72_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07787_ _10017_/A0 _10701_/Q _07817_/S vssd1 vssd1 vccd1 vccd1 _07788_/B sky130_fd_sc_hd__mux2_1
X_09526_ _09529_/A _09526_/B _09526_/C vssd1 vssd1 vccd1 vccd1 _11618_/D sky130_fd_sc_hd__and3_1
XFILLER_83_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06738_ _11332_/Q _06738_/A2 _05789_/Y _06737_/X vssd1 vssd1 vccd1 vccd1 _06738_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _09475_/A _09457_/B vssd1 vssd1 vccd1 vccd1 _09457_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06669_ _10527_/Q _06106_/B _06857_/B1 _11711_/Q _06668_/X vssd1 vssd1 vccd1 vccd1
+ _06669_/X sky130_fd_sc_hd__o221a_1
XFILLER_40_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08408_ _08846_/A0 _11045_/Q _08414_/S vssd1 vssd1 vccd1 vccd1 _08409_/B sky130_fd_sc_hd__mux2_1
X_09388_ _10080_/A0 _11555_/Q _09390_/S vssd1 vssd1 vccd1 vccd1 _11555_/D sky130_fd_sc_hd__mux2_1
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08339_ _08492_/A _08339_/B vssd1 vssd1 vccd1 vccd1 _11012_/D sky130_fd_sc_hd__or2_1
XFILLER_126_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11350_ _11607_/CLK _11350_/D vssd1 vssd1 vccd1 vccd1 _11350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10301_ _11776_/CLK _10301_/D vssd1 vssd1 vccd1 vccd1 _10301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11281_ _11284_/CLK _11281_/D vssd1 vssd1 vccd1 vccd1 _11281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10232_ _11702_/CLK _10232_/D vssd1 vssd1 vccd1 vccd1 _10232_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_133_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10163_ _11793_/Q _10159_/X _10162_/X vssd1 vssd1 vccd1 vccd1 _11793_/D sky130_fd_sc_hd__a21o_1
Xfanout1003 _11867_/A vssd1 vssd1 vccd1 vccd1 _05749_/A sky130_fd_sc_hd__buf_6
XFILLER_43_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1014 _07021_/A vssd1 vssd1 vccd1 vccd1 _10128_/A0 sky130_fd_sc_hd__buf_6
XFILLER_0_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1025 _07018_/A vssd1 vssd1 vccd1 vccd1 _10153_/A1 sky130_fd_sc_hd__buf_6
XFILLER_0_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1036 _10021_/A0 vssd1 vssd1 vccd1 vccd1 _10172_/A1 sky130_fd_sc_hd__buf_6
XFILLER_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1047 _10185_/A0 vssd1 vssd1 vccd1 vccd1 _09396_/A0 sky130_fd_sc_hd__buf_4
X_10094_ _11749_/Q _10104_/B vssd1 vssd1 vccd1 vccd1 _10094_/X sky130_fd_sc_hd__or2_1
XFILLER_86_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1058 input111/X vssd1 vssd1 vccd1 vccd1 _07010_/A sky130_fd_sc_hd__buf_12
Xfanout1069 _10142_/A1 vssd1 vssd1 vccd1 vccd1 _10165_/A1 sky130_fd_sc_hd__buf_6
XFILLER_48_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10996_ _11735_/CLK _10996_/D vssd1 vssd1 vccd1 vccd1 _10996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11617_ _11663_/CLK _11617_/D vssd1 vssd1 vccd1 vccd1 _11617_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11548_ _11675_/CLK _11548_/D vssd1 vssd1 vccd1 vccd1 _11548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11479_ _11485_/CLK _11479_/D vssd1 vssd1 vccd1 vccd1 _11479_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_125_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05971_ _11805_/Q _10180_/A _05969_/X _05970_/X vssd1 vssd1 vccd1 vccd1 _05971_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07710_ _10656_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07710_/X sky130_fd_sc_hd__or2_1
XFILLER_22_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08690_ _08875_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _11199_/D sky130_fd_sc_hd__or2_1
X_07641_ _08441_/B2 _10608_/Q _07642_/S vssd1 vssd1 vccd1 vccd1 _10608_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07572_ _07934_/A _07572_/B vssd1 vssd1 vccd1 vccd1 _10569_/D sky130_fd_sc_hd__or2_1
XFILLER_59_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11607_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09311_ _09995_/A1 _09293_/X _09310_/X _09995_/C1 vssd1 vssd1 vccd1 vccd1 _11506_/D
+ sky130_fd_sc_hd__o211a_1
X_06523_ _10525_/Q _09325_/A _09248_/A _10321_/Q vssd1 vssd1 vccd1 vccd1 _06523_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09242_ _07143_/X _09228_/B _09226_/Y _11473_/Q _09192_/A vssd1 vssd1 vccd1 vccd1
+ _11473_/D sky130_fd_sc_hd__a221o_1
X_06454_ _10590_/Q _06454_/A2 _06539_/B1 _10841_/Q _06624_/C1 vssd1 vssd1 vccd1 vccd1
+ _06454_/X sky130_fd_sc_hd__o221a_2
XFILLER_142_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05405_ _11280_/Q _11279_/Q _05416_/S vssd1 vssd1 vccd1 vccd1 _05406_/D sky130_fd_sc_hd__mux2_1
X_09173_ _10178_/A1 _09171_/B _09173_/B1 vssd1 vssd1 vccd1 vccd1 _09173_/X sky130_fd_sc_hd__a21o_1
X_06385_ _10792_/Q _06540_/A2 _06540_/B1 _10906_/Q vssd1 vssd1 vccd1 vccd1 _06385_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08124_ _10888_/Q _08637_/C vssd1 vssd1 vccd1 vccd1 _08124_/X sky130_fd_sc_hd__or2_1
X_05336_ _11092_/Q _11091_/Q _05372_/S vssd1 vssd1 vccd1 vccd1 _05340_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08055_ _09323_/A0 _10853_/Q _08427_/B vssd1 vssd1 vccd1 vccd1 _08056_/B sky130_fd_sc_hd__mux2_1
XFILLER_135_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05267_ _10440_/Q _10439_/Q _05393_/S vssd1 vssd1 vccd1 vccd1 _05269_/C sky130_fd_sc_hd__mux2_1
XFILLER_116_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07006_ _10266_/Q _08326_/B2 _07038_/S vssd1 vssd1 vccd1 vccd1 _10266_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05198_ _05418_/S _11061_/Q vssd1 vssd1 vccd1 vccd1 _05198_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput106 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 input106/X sky130_fd_sc_hd__clkbuf_2
Xinput117 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 input117/X sky130_fd_sc_hd__clkbuf_16
XFILLER_153_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08957_ _08952_/Y _09830_/B _08956_/X _09959_/B vssd1 vssd1 vccd1 vccd1 _09832_/S
+ sky130_fd_sc_hd__a31o_1
XFILLER_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07908_ _07920_/A _07908_/B vssd1 vssd1 vccd1 vccd1 _10771_/D sky130_fd_sc_hd__or2_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08888_ _11301_/Q _08894_/B vssd1 vssd1 vccd1 vccd1 _08888_/X sky130_fd_sc_hd__or2_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07839_ _07141_/A _07839_/A2 _07961_/S _10734_/Q vssd1 vssd1 vccd1 vccd1 _10734_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _11136_/CLK _10850_/D vssd1 vssd1 vccd1 vccd1 _10850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09509_ _09528_/A _09500_/B _09508_/A _11613_/Q vssd1 vssd1 vccd1 vccd1 _09509_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10781_ _11477_/CLK _10781_/D vssd1 vssd1 vccd1 vccd1 _10781_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11402_ _11411_/CLK _11402_/D vssd1 vssd1 vccd1 vccd1 _11402_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_90 _09232_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11333_ _11657_/CLK _11333_/D vssd1 vssd1 vccd1 vccd1 _11333_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11264_ _11268_/CLK _11264_/D vssd1 vssd1 vccd1 vccd1 _11264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10215_ _11629_/CLK _10215_/D vssd1 vssd1 vccd1 vccd1 _10215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11195_ _11319_/CLK _11195_/D vssd1 vssd1 vccd1 vccd1 _11195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10146_ _10185_/A0 _10154_/B _10150_/B1 vssd1 vssd1 vccd1 vccd1 _10146_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10077_ _10113_/A0 _11737_/Q _10082_/S vssd1 vssd1 vccd1 vccd1 _11737_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10979_ _10981_/CLK _10979_/D vssd1 vssd1 vccd1 vccd1 _10979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06170_ _11798_/Q _10159_/A _09293_/A _11504_/Q vssd1 vssd1 vccd1 vccd1 _06170_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05121_ _11180_/Q _11179_/Q _05399_/S vssd1 vssd1 vccd1 vccd1 _05123_/C sky130_fd_sc_hd__mux2_1
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09860_ _11447_/Q _09879_/A2 _09879_/B1 _10712_/Q _09859_/X vssd1 vssd1 vccd1 vccd1
+ _09861_/D sky130_fd_sc_hd__a221o_4
Xfanout807 _06870_/B1 vssd1 vssd1 vccd1 vccd1 _06999_/A sky130_fd_sc_hd__buf_6
XFILLER_98_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout818 _06166_/A2 vssd1 vssd1 vccd1 vccd1 _06735_/B1 sky130_fd_sc_hd__buf_6
XFILLER_98_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout829 _06161_/A2 vssd1 vssd1 vccd1 vccd1 _07692_/A sky130_fd_sc_hd__buf_4
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _11262_/Q _07630_/B _07630_/Y _08811_/B2 vssd1 vssd1 vccd1 vccd1 _11262_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09791_ _05377_/S _09672_/B _09674_/A _11592_/Q vssd1 vssd1 vccd1 vccd1 _09791_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _08970_/A1 _11228_/Q _08742_/S vssd1 vssd1 vccd1 vccd1 _08743_/B sky130_fd_sc_hd__mux2_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05954_ _11795_/Q _10159_/A _09293_/A _11501_/Q vssd1 vssd1 vccd1 vccd1 _05954_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08673_ _11191_/Q _08705_/B vssd1 vssd1 vccd1 vccd1 _08673_/X sky130_fd_sc_hd__or2_1
XFILLER_22_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05885_ _05656_/X _06622_/A2 _05822_/X _06886_/A2 _05884_/X vssd1 vssd1 vccd1 vccd1
+ _10223_/D sky130_fd_sc_hd__a221o_1
XFILLER_93_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07624_ _08819_/A _08459_/S vssd1 vssd1 vccd1 vccd1 _07624_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07555_ _08987_/A1 _10561_/Q _07557_/S vssd1 vssd1 vccd1 vccd1 _07556_/B sky130_fd_sc_hd__mux2_1
XFILLER_81_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06506_ _10931_/Q _06641_/A2 _08469_/B _11083_/Q vssd1 vssd1 vccd1 vccd1 _06506_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07486_ _10522_/Q _07000_/B _07000_/Y _07451_/B vssd1 vssd1 vccd1 vccd1 _10522_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09225_ _11463_/Q _09205_/Y _09209_/Y _07043_/X vssd1 vssd1 vccd1 vccd1 _11463_/D
+ sky130_fd_sc_hd__a22o_1
X_06437_ _10624_/Q _07939_/A _08286_/A _10723_/Q vssd1 vssd1 vccd1 vccd1 _06437_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09156_ _10161_/A1 _09154_/X _09155_/X _09168_/C1 vssd1 vssd1 vccd1 vccd1 _11422_/D
+ sky130_fd_sc_hd__o211a_1
X_06368_ _10704_/Q _06807_/A2 _06728_/B1 _10538_/Q _06367_/X vssd1 vssd1 vccd1 vccd1
+ _06368_/X sky130_fd_sc_hd__o221a_1
XFILLER_147_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08107_ _08819_/A _08107_/B vssd1 vssd1 vccd1 vccd1 _10878_/D sky130_fd_sc_hd__or2_1
X_05319_ _10608_/Q _10607_/Q _05391_/S vssd1 vssd1 vccd1 vccd1 _05323_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09087_ _09276_/A1 _09099_/B _08873_/A vssd1 vssd1 vccd1 vccd1 _09087_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06299_ _06296_/X _06298_/X _07297_/A _06294_/X vssd1 vssd1 vccd1 vccd1 _06299_/X
+ sky130_fd_sc_hd__a211o_1
X_08038_ _08853_/A1 _08035_/S _08037_/X _08843_/C1 vssd1 vssd1 vccd1 vccd1 _10843_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10000_ _10110_/A0 _11687_/Q _10008_/S vssd1 vssd1 vccd1 vccd1 _11687_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09989_ _11681_/Q _09977_/X _09988_/X vssd1 vssd1 vccd1 vccd1 _11681_/D sky130_fd_sc_hd__a21o_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10902_ _11280_/CLK _10902_/D vssd1 vssd1 vccd1 vccd1 _10902_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10833_ _11601_/CLK _10833_/D vssd1 vssd1 vccd1 vccd1 _10833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10764_ _10769_/CLK _10764_/D vssd1 vssd1 vccd1 vccd1 _10764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10695_ _11744_/CLK _10695_/D vssd1 vssd1 vccd1 vccd1 _10695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11316_ _11385_/CLK _11316_/D vssd1 vssd1 vccd1 vccd1 _11316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11247_ _11251_/CLK _11247_/D vssd1 vssd1 vccd1 vccd1 _11247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11178_ _11268_/CLK _11178_/D vssd1 vssd1 vccd1 vccd1 _11178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10129_ _07057_/A _11775_/Q _10135_/S vssd1 vssd1 vccd1 vccd1 _11775_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05670_ _11191_/Q _05531_/Y _05555_/Y _11200_/Q vssd1 vssd1 vccd1 vccd1 _05679_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07340_ _10436_/Q _07350_/S _07346_/B1 _07005_/A vssd1 vssd1 vccd1 vccd1 _10436_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_143_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07271_ _08789_/A1 _10404_/Q _09187_/S vssd1 vssd1 vccd1 vccd1 _07272_/B sky130_fd_sc_hd__mux2_1
XFILLER_91_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09010_ _10153_/A1 _08994_/X _09009_/X _09032_/C1 vssd1 vssd1 vccd1 vccd1 _11356_/D
+ sky130_fd_sc_hd__o211a_1
X_06222_ _11429_/Q _09154_/A _06221_/X _06357_/C1 vssd1 vssd1 vccd1 vccd1 _06222_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06153_ _11772_/Q _05865_/B _08647_/B _10303_/Q _06152_/X vssd1 vssd1 vccd1 vccd1
+ _06153_/X sky130_fd_sc_hd__o221a_1
XFILLER_145_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05104_ _11262_/Q _11261_/Q _05392_/S vssd1 vssd1 vccd1 vccd1 _05107_/B sky130_fd_sc_hd__mux2_1
X_06084_ _11751_/Q _10087_/A _10137_/A _11787_/Q _06349_/C1 vssd1 vssd1 vccd1 vccd1
+ _06084_/X sky130_fd_sc_hd__o221a_1
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09912_ _10363_/Q _09572_/A _09565_/B _10356_/Q _09911_/X vssd1 vssd1 vccd1 vccd1
+ _09917_/B sky130_fd_sc_hd__a221o_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout604 _06430_/A2 vssd1 vssd1 vccd1 vccd1 _06643_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_67_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout615 _05737_/X vssd1 vssd1 vccd1 vccd1 _07300_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_154_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout626 _05737_/X vssd1 vssd1 vccd1 vccd1 _06696_/A2 sky130_fd_sc_hd__buf_4
XFILLER_113_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _10781_/Q _09883_/B1 _09881_/B1 _10772_/Q vssd1 vssd1 vccd1 vccd1 _09843_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout637 _05100_/Y vssd1 vssd1 vccd1 vccd1 _09447_/B sky130_fd_sc_hd__buf_8
XFILLER_99_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout648 _05072_/Y vssd1 vssd1 vccd1 vccd1 _09525_/A sky130_fd_sc_hd__buf_4
XFILLER_150_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout659 _11627_/Q vssd1 vssd1 vccd1 vccd1 _05626_/A2 sky130_fd_sc_hd__clkbuf_16
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _10185_/A0 _06976_/X _06985_/X _06996_/C1 vssd1 vssd1 vccd1 vccd1 _10260_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _11650_/Q _11649_/Q _11648_/Q _11647_/Q vssd1 vssd1 vccd1 vccd1 _09775_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ _08810_/A _08725_/B vssd1 vssd1 vccd1 vccd1 _11219_/D sky130_fd_sc_hd__or2_1
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05937_ _10835_/Q _06539_/B1 _06455_/B1 _10428_/Q _05936_/X vssd1 vssd1 vccd1 vccd1
+ _05937_/X sky130_fd_sc_hd__o221a_2
XFILLER_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _08092_/X _08742_/S _08655_/X _08427_/A vssd1 vssd1 vccd1 vccd1 _11183_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05868_ _10602_/Q _06635_/B1 _06556_/B1 _11175_/Q _05867_/X vssd1 vssd1 vccd1 vccd1
+ _05868_/X sky130_fd_sc_hd__o221a_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _10587_/Q _07597_/Y _07600_/Y _07022_/X vssd1 vssd1 vccd1 vccd1 _10587_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _11149_/Q _08591_/B vssd1 vssd1 vccd1 vccd1 _08587_/X sky130_fd_sc_hd__or2_1
X_05799_ _10455_/Q _06643_/A2 _10119_/A _10451_/Q vssd1 vssd1 vccd1 vccd1 _05799_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_23_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07538_ _07042_/A _07513_/S _07537_/X _07868_/C1 vssd1 vssd1 vccd1 vccd1 _10553_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07469_ _08931_/A1 _10512_/Q _07477_/S vssd1 vssd1 vccd1 vccd1 _07470_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09208_ _09228_/A _09208_/B vssd1 vssd1 vccd1 vccd1 _09208_/Y sky130_fd_sc_hd__nor2_2
XFILLER_155_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10480_ _11719_/CLK _10480_/D vssd1 vssd1 vccd1 vccd1 _10480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09139_ _11415_/Q _09149_/B vssd1 vssd1 vccd1 vccd1 _09139_/X sky130_fd_sc_hd__or2_1
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11101_ _11186_/CLK _11101_/D vssd1 vssd1 vccd1 vccd1 _11101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11032_ _11607_/CLK _11032_/D vssd1 vssd1 vccd1 vccd1 _11032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_wb_clk_i clkbuf_4_10__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10782_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10816_ _11641_/CLK _10816_/D vssd1 vssd1 vccd1 vccd1 _10816_/Q sky130_fd_sc_hd__dfxtp_1
X_11796_ _11801_/CLK _11796_/D vssd1 vssd1 vccd1 vccd1 _11796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10747_ _10804_/CLK _10747_/D vssd1 vssd1 vccd1 vccd1 _10747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10678_ _11471_/CLK _10678_/D vssd1 vssd1 vccd1 vccd1 _10678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput207 _05482_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_4
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06840_ _11334_/Q _06704_/B _06839_/X vssd1 vssd1 vccd1 vccd1 _10248_/D sky130_fd_sc_hd__a21o_1
XFILLER_110_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06771_ _10694_/Q _07203_/A _06858_/B1 _10518_/Q vssd1 vssd1 vccd1 vccd1 _06771_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08510_ _09275_/A1 _08529_/S _08509_/X _09092_/C1 vssd1 vssd1 vccd1 vccd1 _11104_/D
+ sky130_fd_sc_hd__o211a_1
X_05722_ _10961_/Q _05537_/Y _05573_/Y _10964_/Q _05721_/X vssd1 vssd1 vccd1 vccd1
+ _05728_/B sky130_fd_sc_hd__a221o_1
XFILLER_97_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09490_ _09490_/A vssd1 vssd1 vccd1 vccd1 _09490_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08441_ _11062_/Q _08437_/Y _08438_/Y _08441_/B2 vssd1 vssd1 vccd1 vccd1 _11062_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05653_ _11293_/Q _05549_/Y _05650_/X _05652_/X vssd1 vssd1 vccd1 vccd1 _05653_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_36_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08372_ _10149_/A1 _11028_/Q _08439_/B vssd1 vssd1 vccd1 vccd1 _08373_/B sky130_fd_sc_hd__mux2_1
X_05584_ _05076_/A _11385_/Q _11380_/Q _05620_/B2 _05583_/X vssd1 vssd1 vccd1 vccd1
+ _05585_/B sky130_fd_sc_hd__a221o_4
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07323_ _09206_/A _08162_/S vssd1 vssd1 vccd1 vccd1 _07323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07254_ _07254_/A _07854_/B vssd1 vssd1 vccd1 vccd1 _07259_/S sky130_fd_sc_hd__or2_4
XFILLER_137_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06205_ _11245_/Q _08765_/A _06201_/X _06204_/X vssd1 vssd1 vccd1 vccd1 _06205_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07185_ _07141_/A _07172_/S _07184_/X _07884_/C1 vssd1 vssd1 vccd1 vccd1 _10353_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06136_ _10647_/Q _07692_/A _06132_/X _06135_/X vssd1 vssd1 vccd1 vccd1 _06136_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06067_ _11279_/Q _06454_/A2 _06455_/B1 _10429_/Q _06066_/X vssd1 vssd1 vccd1 vccd1
+ _06067_/X sky130_fd_sc_hd__o221a_2
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout401 _05423_/Y vssd1 vssd1 vccd1 vccd1 _09881_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_99_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout412 _05357_/Y vssd1 vssd1 vccd1 vccd1 _09570_/B sky130_fd_sc_hd__buf_8
Xfanout423 _05302_/Y vssd1 vssd1 vccd1 vccd1 _09871_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout434 _05238_/X vssd1 vssd1 vccd1 vccd1 _09568_/D sky130_fd_sc_hd__buf_8
XFILLER_101_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout445 _05179_/Y vssd1 vssd1 vccd1 vccd1 _09881_/A2 sky130_fd_sc_hd__buf_4
XFILLER_59_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout456 _05113_/Y vssd1 vssd1 vccd1 vccd1 _09571_/A sky130_fd_sc_hd__buf_8
X_09826_ _09561_/B _09823_/B _09600_/B vssd1 vssd1 vccd1 vccd1 _09827_/B sky130_fd_sc_hd__o21ba_1
Xfanout467 _09022_/C1 vssd1 vssd1 vccd1 vccd1 _08588_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout478 _06899_/X vssd1 vssd1 vccd1 vccd1 _07018_/B sky130_fd_sc_hd__buf_6
Xfanout489 fanout510/X vssd1 vssd1 vccd1 vccd1 _07882_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09757_ _09757_/A _09757_/B _09757_/C _09757_/D vssd1 vssd1 vccd1 vccd1 _09758_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_74_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _10929_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_06969_ _09539_/B _06968_/X _06969_/S vssd1 vssd1 vccd1 vccd1 _06969_/X sky130_fd_sc_hd__mux2_4
XFILLER_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _08875_/A _08708_/B vssd1 vssd1 vccd1 vccd1 _11208_/D sky130_fd_sc_hd__or2_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09688_ _09703_/A _09688_/B vssd1 vssd1 vccd1 vccd1 _11636_/D sky130_fd_sc_hd__or2_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _11174_/Q _08437_/A _08146_/S _08438_/A vssd1 vssd1 vccd1 vccd1 _08639_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11650_/CLK _11650_/D vssd1 vssd1 vccd1 vccd1 _11650_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10601_ _11262_/CLK _10601_/D vssd1 vssd1 vccd1 vccd1 _10601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11581_ _11584_/CLK _11581_/D vssd1 vssd1 vccd1 vccd1 _11581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10532_ _11745_/CLK _10532_/D vssd1 vssd1 vccd1 vccd1 _10532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10463_ _11136_/CLK _10463_/D vssd1 vssd1 vccd1 vccd1 _10463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10394_ _10735_/CLK _10394_/D vssd1 vssd1 vccd1 vccd1 _10394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11015_ _11023_/CLK _11015_/D vssd1 vssd1 vccd1 vccd1 _11015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout990 _11869_/A vssd1 vssd1 vccd1 vccd1 _06550_/C1 sky130_fd_sc_hd__buf_6
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1081 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1081/HI io_oeb[11] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_1092 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1092/HI io_oeb[22] sky130_fd_sc_hd__conb_1
XFILLER_127_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11779_ _11779_/CLK _11779_/D vssd1 vssd1 vccd1 vccd1 _11779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_75_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11291_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08990_ _09172_/A1 _08972_/X _08989_/X _09122_/C1 vssd1 vssd1 vccd1 vccd1 _11347_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07941_ _08902_/B _08085_/B vssd1 vssd1 vccd1 vccd1 _07941_/Y sky130_fd_sc_hd__nor2_2
XFILLER_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07872_ _08684_/A _07872_/B vssd1 vssd1 vccd1 vccd1 _10754_/D sky130_fd_sc_hd__or2_1
XFILLER_96_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09611_ _10631_/Q _09909_/A2 _09573_/C _10392_/Q _09604_/X vssd1 vssd1 vccd1 vccd1
+ _09615_/A sky130_fd_sc_hd__a221o_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06823_ _06813_/X _06814_/X _06817_/X _06822_/X vssd1 vssd1 vccd1 vccd1 _06823_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06754_ _06853_/A1 _10242_/Q _06852_/A3 _06743_/X _06753_/X vssd1 vssd1 vccd1 vccd1
+ _06754_/X sky130_fd_sc_hd__a32o_1
X_09542_ _09539_/X _09661_/B _09959_/B vssd1 vssd1 vccd1 vccd1 _09542_/X sky130_fd_sc_hd__a21o_2
XFILLER_110_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05705_ _11050_/Q _05543_/Y _05615_/Y _11046_/Q vssd1 vssd1 vccd1 vccd1 _05709_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06685_ _11712_/Q _06685_/B vssd1 vssd1 vccd1 vccd1 _06685_/X sky130_fd_sc_hd__or2_1
X_09473_ _09441_/B input16/X _09441_/Y input34/X _09472_/X vssd1 vssd1 vccd1 vccd1
+ _09473_/X sky130_fd_sc_hd__a221o_1
XFILLER_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08424_ _08902_/B _08426_/B vssd1 vssd1 vccd1 vccd1 _08424_/Y sky130_fd_sc_hd__nor2_2
X_05636_ _11319_/Q _05537_/Y _05573_/Y _11322_/Q _05525_/X vssd1 vssd1 vccd1 vccd1
+ _05644_/B sky130_fd_sc_hd__a221o_1
XFILLER_52_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08355_ _08492_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _11020_/D sky130_fd_sc_hd__or2_1
X_05567_ _05567_/A _05567_/B vssd1 vssd1 vccd1 vccd1 _05567_/Y sky130_fd_sc_hd__nor2_8
XFILLER_138_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07306_ _08439_/A _08760_/S vssd1 vssd1 vccd1 vccd1 _07306_/Y sky130_fd_sc_hd__nand2_2
X_08286_ _08286_/A _08649_/B _08649_/C vssd1 vssd1 vccd1 vccd1 _08467_/S sky130_fd_sc_hd__and3_4
XFILLER_138_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05498_ _10243_/Q input55/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05498_/X sky130_fd_sc_hd__mux2_1
X_07237_ _08647_/A _07663_/S _07420_/A vssd1 vssd1 vccd1 vccd1 _07237_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07168_ _08929_/A1 _10345_/Q _07172_/S vssd1 vssd1 vccd1 vccd1 _07169_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06119_ _06119_/A _06119_/B _06119_/C vssd1 vssd1 vccd1 vccd1 _06119_/X sky130_fd_sc_hd__and3_2
XFILLER_156_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07099_ _10305_/Q _07098_/X _07109_/S vssd1 vssd1 vccd1 vccd1 _10305_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout220 _07346_/B1 vssd1 vssd1 vccd1 vccd1 _07846_/S sky130_fd_sc_hd__buf_6
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout231 _07491_/S vssd1 vssd1 vccd1 vccd1 _07490_/S sky130_fd_sc_hd__buf_6
XFILLER_8_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout242 _09488_/Y vssd1 vssd1 vccd1 vccd1 _09489_/C sky130_fd_sc_hd__buf_4
Xfanout253 _08707_/S vssd1 vssd1 vccd1 vccd1 _08695_/S sky130_fd_sc_hd__buf_6
Xfanout264 _08404_/S vssd1 vssd1 vccd1 vccd1 _08414_/S sky130_fd_sc_hd__buf_6
Xfanout275 _08123_/X vssd1 vssd1 vccd1 vccd1 _08146_/S sky130_fd_sc_hd__buf_4
Xfanout286 _07854_/X vssd1 vssd1 vccd1 vccd1 _07890_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09809_ _10299_/Q _09909_/A2 _09953_/B1 _10532_/Q _09804_/X vssd1 vssd1 vccd1 vccd1
+ _09811_/C sky130_fd_sc_hd__a221o_2
Xfanout297 _08102_/S vssd1 vssd1 vccd1 vccd1 _08120_/S sky130_fd_sc_hd__buf_6
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _11702_/CLK _11702_/D vssd1 vssd1 vccd1 vccd1 _11702_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11633_/CLK _11633_/D vssd1 vssd1 vccd1 vccd1 _11633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11564_ _11763_/CLK _11564_/D vssd1 vssd1 vccd1 vccd1 _11564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10515_ _10735_/CLK _10515_/D vssd1 vssd1 vccd1 vccd1 _10515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11495_ _11495_/CLK _11495_/D vssd1 vssd1 vccd1 vccd1 _11495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10446_ _11780_/CLK _10446_/D vssd1 vssd1 vccd1 vccd1 _10446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _11474_/CLK _10377_/D vssd1 vssd1 vccd1 vccd1 _10377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_122_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11711_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06470_ _11228_/Q _06470_/A2 _06640_/B1 _11310_/Q vssd1 vssd1 vccd1 vccd1 _06470_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 _10086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_191 _07059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05421_ _10424_/Q _10423_/Q _06945_/B vssd1 vssd1 vccd1 vccd1 _05422_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08140_ _08970_/A1 _10896_/Q _08140_/S vssd1 vssd1 vccd1 vccd1 _08141_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05352_ _11140_/Q _11139_/Q _05377_/S vssd1 vssd1 vccd1 vccd1 _05354_/C sky130_fd_sc_hd__mux2_2
XFILLER_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08071_ _10861_/Q _08085_/B vssd1 vssd1 vccd1 vccd1 _08071_/X sky130_fd_sc_hd__or2_1
XFILLER_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05283_ _05426_/S _11173_/Q _10894_/Q _09681_/A _05282_/X vssd1 vssd1 vccd1 vccd1
+ _05291_/A sky130_fd_sc_hd__a221o_2
XFILLER_88_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07022_ _07333_/A _07022_/B vssd1 vssd1 vccd1 vccd1 _07022_/X sky130_fd_sc_hd__or2_4
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08973_ _11339_/Q _08989_/B vssd1 vssd1 vccd1 vccd1 _08973_/X sky130_fd_sc_hd__or2_1
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07924_ _07934_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _10779_/D sky130_fd_sc_hd__or2_1
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07855_ _10746_/Q _07893_/B vssd1 vssd1 vccd1 vccd1 _07855_/X sky130_fd_sc_hd__or2_1
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06806_ _10578_/Q _06806_/A2 _06806_/B1 _10677_/Q vssd1 vssd1 vccd1 vccd1 _06806_/X
+ sky130_fd_sc_hd__o22a_1
X_07786_ _07928_/A _07786_/B vssd1 vssd1 vccd1 vccd1 _10700_/D sky130_fd_sc_hd__or2_1
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ _09525_/A _09528_/B _09495_/C vssd1 vssd1 vccd1 vccd1 _09526_/C sky130_fd_sc_hd__or3b_1
XFILLER_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06737_ _11122_/Q _06737_/A2 _06737_/B1 _10974_/Q _06736_/X vssd1 vssd1 vccd1 vccd1
+ _06737_/X sky130_fd_sc_hd__o221a_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_06668_ _10370_/Q _06799_/A2 _06871_/B1 _10729_/Q vssd1 vssd1 vccd1 vccd1 _06668_/X
+ sky130_fd_sc_hd__o22a_1
X_09456_ input35/X _09442_/X _09455_/X vssd1 vssd1 vccd1 vccd1 _09457_/B sky130_fd_sc_hd__o21ai_1
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05619_ _05619_/A1 _11378_/Q _11374_/Q _05619_/B2 _05617_/X vssd1 vssd1 vccd1 vccd1
+ _05619_/X sky130_fd_sc_hd__a221o_1
X_08407_ _08851_/A _08407_/B vssd1 vssd1 vccd1 vccd1 _11044_/D sky130_fd_sc_hd__or2_1
XFILLER_61_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09387_ _10115_/A0 _11554_/Q _09390_/S vssd1 vssd1 vccd1 vccd1 _11554_/D sky130_fd_sc_hd__mux2_1
X_06599_ _10472_/Q _06642_/A2 _06598_/X _06642_/C1 vssd1 vssd1 vccd1 vccd1 _06599_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08338_ _09393_/A0 _11012_/Q _08360_/S vssd1 vssd1 vccd1 vccd1 _08339_/B sky130_fd_sc_hd__mux2_1
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08269_ _08771_/A _08269_/B vssd1 vssd1 vccd1 vccd1 _10966_/D sky130_fd_sc_hd__or2_1
XFILLER_119_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10300_ _11766_/CLK _10300_/D vssd1 vssd1 vccd1 vccd1 _10300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11280_ _11280_/CLK _11280_/D vssd1 vssd1 vccd1 vccd1 _11280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10231_ _11665_/CLK _10231_/D vssd1 vssd1 vccd1 vccd1 _10231_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10162_ _10162_/A1 _10176_/B _10166_/B1 vssd1 vssd1 vccd1 vccd1 _10162_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1004 input80/X vssd1 vssd1 vccd1 vccd1 _11867_/A sky130_fd_sc_hd__buf_4
Xfanout1015 _10105_/A1 vssd1 vssd1 vccd1 vccd1 _09323_/A0 sky130_fd_sc_hd__buf_4
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1026 input115/X vssd1 vssd1 vccd1 vccd1 _07018_/A sky130_fd_sc_hd__buf_12
X_10093_ _11748_/Q _10087_/X _10092_/X vssd1 vssd1 vccd1 vccd1 _11748_/D sky130_fd_sc_hd__a21o_1
Xfanout1037 input114/X vssd1 vssd1 vccd1 vccd1 _10021_/A0 sky130_fd_sc_hd__buf_12
Xfanout1048 _07092_/A vssd1 vssd1 vccd1 vccd1 _10185_/A0 sky130_fd_sc_hd__buf_6
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1059 _10166_/A1 vssd1 vssd1 vccd1 vccd1 _09985_/A1 sky130_fd_sc_hd__buf_6
XFILLER_134_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10995_ _11735_/CLK _10995_/D vssd1 vssd1 vccd1 vccd1 _10995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11616_ _11812_/CLK _11616_/D vssd1 vssd1 vccd1 vccd1 _11616_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ _11791_/CLK _11547_/D vssd1 vssd1 vccd1 vccd1 _11547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11478_ _11485_/CLK _11478_/D vssd1 vssd1 vccd1 vccd1 _11478_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10429_ _11280_/CLK _10429_/D vssd1 vssd1 vccd1 vccd1 _10429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05970_ _10259_/Q _06230_/A2 _06903_/A _10196_/Q vssd1 vssd1 vccd1 vccd1 _05970_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_61_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07640_ _08440_/B2 _10607_/Q _07642_/S vssd1 vssd1 vccd1 vccd1 _10607_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07571_ _07211_/A _10569_/Q _07591_/S vssd1 vssd1 vccd1 vccd1 _07572_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09310_ _11506_/Q _09310_/B vssd1 vssd1 vccd1 vccd1 _09310_/X sky130_fd_sc_hd__or2_1
X_06522_ _10626_/Q _07939_/A _08286_/A _10725_/Q vssd1 vssd1 vccd1 vccd1 _06522_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09241_ _09226_/A _09240_/X _09241_/B1 vssd1 vssd1 vccd1 vccd1 _11472_/D sky130_fd_sc_hd__o21a_1
XFILLER_61_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06453_ _11066_/Q _06538_/A2 _06453_/B1 _10644_/Q vssd1 vssd1 vccd1 vccd1 _06453_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_90_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11661_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_05404_ _10584_/Q _10583_/Q _06939_/A vssd1 vssd1 vccd1 vccd1 _05406_/C sky130_fd_sc_hd__mux2_1
X_09172_ _09172_/A1 _09154_/X _09171_/X _10175_/C1 vssd1 vssd1 vccd1 vccd1 _11430_/D
+ sky130_fd_sc_hd__o211a_1
X_06384_ _10588_/Q _06454_/A2 _06539_/B1 _10839_/Q _06624_/C1 vssd1 vssd1 vccd1 vccd1
+ _06387_/B sky130_fd_sc_hd__o221a_1
X_08123_ _08123_/A _10119_/B _09038_/C vssd1 vssd1 vccd1 vccd1 _08123_/X sky130_fd_sc_hd__or3_1
X_05335_ _05335_/A _05335_/B vssd1 vssd1 vccd1 vccd1 _05335_/Y sky130_fd_sc_hd__nor2_8
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08054_ _08054_/A _10119_/B _09038_/C vssd1 vssd1 vccd1 vccd1 _08427_/B sky130_fd_sc_hd__or3_4
X_05266_ _10443_/Q _10738_/Q _05394_/S vssd1 vssd1 vccd1 vccd1 _05269_/B sky130_fd_sc_hd__mux2_1
X_07005_ _07005_/A _07599_/A vssd1 vssd1 vccd1 vccd1 _07005_/X sky130_fd_sc_hd__or2_4
XFILLER_66_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05197_ _05418_/S _11062_/Q vssd1 vssd1 vccd1 vccd1 _05197_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_103_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput107 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 _07147_/A sky130_fd_sc_hd__buf_4
Xinput118 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _05729_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08956_ _09538_/A _08956_/B _11587_/Q _09491_/C vssd1 vssd1 vccd1 vccd1 _08956_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_5_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07907_ _10019_/A0 _10771_/Q _09221_/C vssd1 vssd1 vccd1 vccd1 _07908_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08887_ _08941_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _11300_/D sky130_fd_sc_hd__or2_1
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07838_ _10051_/A1 _07839_/A2 _07961_/S _10733_/Q vssd1 vssd1 vccd1 vccd1 _10733_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07769_ _10689_/Q _07316_/X _07773_/S vssd1 vssd1 vccd1 vccd1 _10689_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09508_ _09508_/A vssd1 vssd1 vccd1 vccd1 _09508_/Y sky130_fd_sc_hd__inv_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10780_ _11470_/CLK _10780_/D vssd1 vssd1 vccd1 vccd1 _10780_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _11592_/Q _11651_/Q _09440_/S vssd1 vssd1 vccd1 vccd1 _11592_/D sky130_fd_sc_hd__mux2_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11401_ _11745_/CLK _11401_/D vssd1 vssd1 vccd1 vccd1 _11401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_80 _11623_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_91 _09229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11332_ _11332_/CLK _11332_/D vssd1 vssd1 vccd1 vccd1 _11332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11263_ _11268_/CLK _11263_/D vssd1 vssd1 vccd1 vccd1 _11263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10214_ _11629_/CLK _10214_/D vssd1 vssd1 vccd1 vccd1 _10214_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11194_ _11325_/CLK _11194_/D vssd1 vssd1 vccd1 vccd1 _11194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10145_ _10184_/A0 _10137_/X _10144_/X _10155_/C1 vssd1 vssd1 vccd1 vccd1 _11785_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10076_ _10112_/A0 _11736_/Q _10082_/S vssd1 vssd1 vccd1 vccd1 _11736_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10978_ _11224_/CLK _10978_/D vssd1 vssd1 vccd1 vccd1 _10978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05120_ _10309_/Q _10308_/Q _06942_/B vssd1 vssd1 vccd1 vccd1 _05123_/B sky130_fd_sc_hd__mux2_1
XFILLER_15_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout808 _06166_/A2 vssd1 vssd1 vccd1 vccd1 _06870_/B1 sky130_fd_sc_hd__buf_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout819 _05745_/X vssd1 vssd1 vccd1 vccd1 _06166_/A2 sky130_fd_sc_hd__buf_12
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _08810_/A _08810_/B vssd1 vssd1 vccd1 vccd1 _11261_/D sky130_fd_sc_hd__or2_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _11650_/Q _08950_/B _09789_/X _09407_/A vssd1 vssd1 vccd1 vccd1 _11650_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _08969_/A1 _08748_/S _08740_/X _08821_/A vssd1 vssd1 vccd1 vccd1 _11227_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05953_ _11749_/Q _05953_/A2 _08994_/A _11785_/Q _06349_/C1 vssd1 vssd1 vccd1 vccd1
+ _05953_/X sky130_fd_sc_hd__o221a_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08672_ _08873_/A _08672_/B vssd1 vssd1 vccd1 vccd1 _11190_/D sky130_fd_sc_hd__or2_1
X_05884_ _06535_/A _05822_/X _05883_/X _06664_/C1 vssd1 vssd1 vccd1 vccd1 _05884_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07623_ _09976_/A _08560_/C _07847_/C vssd1 vssd1 vccd1 vccd1 _07623_/X sky130_fd_sc_hd__and3_2
XFILLER_148_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07554_ _07926_/A _07554_/B vssd1 vssd1 vccd1 vccd1 _10560_/D sky130_fd_sc_hd__or2_1
XFILLER_59_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06505_ _06501_/X _06502_/X _06504_/X _07689_/A vssd1 vssd1 vccd1 vccd1 _06505_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07485_ _10521_/Q _07000_/B _07000_/Y _07143_/X vssd1 vssd1 vccd1 vccd1 _10521_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09224_ _11462_/Q _09205_/Y _09209_/Y _07040_/X vssd1 vssd1 vccd1 vccd1 _11462_/D
+ sky130_fd_sc_hd__a22o_1
X_06436_ _10774_/Q _06646_/A2 _06432_/X _06435_/X vssd1 vssd1 vccd1 vccd1 _06436_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_107_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09155_ _11422_/Q _09171_/B vssd1 vssd1 vccd1 vccd1 _09155_/X sky130_fd_sc_hd__or2_1
X_06367_ _10773_/Q _06862_/A2 _06806_/B1 _10662_/Q vssd1 vssd1 vccd1 vccd1 _06367_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08106_ _10878_/Q _07052_/A _08120_/S vssd1 vssd1 vccd1 vccd1 _08107_/B sky130_fd_sc_hd__mux2_1
X_05318_ _05318_/A _05318_/B _05318_/C _05318_/D vssd1 vssd1 vccd1 vccd1 _05324_/A
+ sky130_fd_sc_hd__or4_4
X_06298_ _11754_/Q _06413_/A2 _06363_/A2 _11486_/Q _06297_/X vssd1 vssd1 vccd1 vccd1
+ _06298_/X sky130_fd_sc_hd__o221a_1
X_09086_ _11390_/Q _09082_/X _09085_/X vssd1 vssd1 vccd1 vccd1 _11390_/D sky130_fd_sc_hd__a21o_1
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05249_ _10976_/Q _10975_/Q _05380_/S vssd1 vssd1 vccd1 vccd1 _05253_/A sky130_fd_sc_hd__mux2_1
X_08037_ _10843_/Q _08037_/B vssd1 vssd1 vccd1 vccd1 _08037_/X sky130_fd_sc_hd__or2_1
XFILLER_122_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09988_ _10171_/A1 _09994_/B _10178_/B1 vssd1 vssd1 vccd1 vccd1 _09988_/X sky130_fd_sc_hd__a21o_1
XFILLER_104_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08939_ _08939_/A1 _08940_/S _08938_/X _08943_/C1 vssd1 vssd1 vccd1 vccd1 _11328_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ _11005_/CLK _10901_/D vssd1 vssd1 vccd1 vccd1 _10901_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10832_ _11151_/CLK _10832_/D vssd1 vssd1 vccd1 vccd1 _10832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10763_ _11458_/CLK _10763_/D vssd1 vssd1 vccd1 vccd1 _10763_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_13_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ _11719_/CLK _10694_/D vssd1 vssd1 vccd1 vccd1 _10694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11315_ _11385_/CLK _11315_/D vssd1 vssd1 vccd1 vccd1 _11315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11246_ _11575_/CLK _11246_/D vssd1 vssd1 vccd1 vccd1 _11246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11177_ _11177_/CLK _11177_/D vssd1 vssd1 vccd1 vccd1 _11177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10128_ _10128_/A0 _11774_/Q _10135_/S vssd1 vssd1 vccd1 vccd1 _11774_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10059_ _11721_/Q _10028_/B _10085_/S _07037_/B vssd1 vssd1 vccd1 vccd1 _11721_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11601_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07270_ _07796_/A _07270_/B vssd1 vssd1 vccd1 vccd1 _10403_/D sky130_fd_sc_hd__or2_1
XFILLER_108_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06221_ _11376_/Q _06221_/A2 _09110_/A _11409_/Q _06220_/X vssd1 vssd1 vccd1 vccd1
+ _06221_/X sky130_fd_sc_hd__o221a_2
XFILLER_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06152_ _11075_/Q _06152_/B vssd1 vssd1 vccd1 vccd1 _06152_/X sky130_fd_sc_hd__or2_1
XFILLER_144_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05103_ _10602_/Q _10601_/Q _05391_/S vssd1 vssd1 vccd1 vccd1 _05107_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06083_ _11523_/Q _09326_/A _06363_/A2 _11483_/Q vssd1 vssd1 vccd1 vccd1 _06083_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09911_ _10481_/Q _09571_/B _09567_/B _10489_/Q vssd1 vssd1 vccd1 vccd1 _09911_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout605 _06430_/A2 vssd1 vssd1 vccd1 vccd1 _07046_/A sky130_fd_sc_hd__buf_8
Xfanout616 _06748_/A2 vssd1 vssd1 vccd1 vccd1 _06873_/A2 sky130_fd_sc_hd__buf_6
XFILLER_99_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout627 _05736_/Y vssd1 vssd1 vccd1 vccd1 _09059_/A sky130_fd_sc_hd__clkbuf_16
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _09842_/A _09842_/B _09842_/C _09842_/D vssd1 vssd1 vccd1 vccd1 _09850_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_59_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout638 _05079_/Y vssd1 vssd1 vccd1 vccd1 _05630_/B1 sky130_fd_sc_hd__clkbuf_16
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout649 _05072_/Y vssd1 vssd1 vccd1 vccd1 _09528_/A sky130_fd_sc_hd__buf_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _11647_/Q _09771_/Y _09772_/X _09554_/B _09406_/B vssd1 vssd1 vccd1 vccd1
+ _09773_/X sky130_fd_sc_hd__o221a_1
X_06985_ _10260_/Q _06995_/B vssd1 vssd1 vccd1 vccd1 _06985_/X sky130_fd_sc_hd__or2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08724_ _11219_/Q _08818_/A1 _08726_/S vssd1 vssd1 vccd1 vccd1 _08725_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05936_ _10583_/Q _06454_/A2 _06455_/A2 _10862_/Q vssd1 vssd1 vccd1 vccd1 _05936_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_113_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08655_ _11183_/Q _08655_/B _08750_/B vssd1 vssd1 vccd1 vccd1 _08655_/X sky130_fd_sc_hd__or3_1
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05867_ _11070_/Q _06731_/B1 _06637_/A2 _10743_/Q vssd1 vssd1 vccd1 vccd1 _05867_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _10586_/Q _07598_/Y _07599_/Y _07232_/X vssd1 vssd1 vccd1 vccd1 _10586_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _08757_/A _08586_/B vssd1 vssd1 vccd1 vccd1 _11148_/D sky130_fd_sc_hd__or2_1
X_05798_ _10909_/Q _07046_/A _05794_/X _05797_/X vssd1 vssd1 vccd1 vccd1 _05798_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07537_ _10553_/Q _07537_/B vssd1 vssd1 vccd1 vccd1 _07537_/X sky130_fd_sc_hd__or2_1
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07468_ _07476_/A _07468_/B vssd1 vssd1 vccd1 vccd1 _10511_/D sky130_fd_sc_hd__or2_1
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ _07303_/X _09221_/C _09206_/Y _11451_/Q _09229_/A vssd1 vssd1 vccd1 vccd1
+ _11451_/D sky130_fd_sc_hd__o221a_1
X_06419_ _10895_/Q _08123_/A _06415_/X _06418_/X vssd1 vssd1 vccd1 vccd1 _06420_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_120_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07399_ _10015_/A0 _10476_/Q _07437_/S vssd1 vssd1 vccd1 vccd1 _07400_/B sky130_fd_sc_hd__mux2_1
XFILLER_120_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09138_ _11414_/Q _09132_/X _09137_/X vssd1 vssd1 vccd1 vccd1 _11414_/D sky130_fd_sc_hd__a21o_1
XFILLER_147_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09069_ _11383_/Q _09077_/B vssd1 vssd1 vccd1 vccd1 _09069_/X sky130_fd_sc_hd__or2_1
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11100_ _11186_/CLK _11100_/D vssd1 vssd1 vccd1 vccd1 _11100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11031_ _11607_/CLK _11031_/D vssd1 vssd1 vccd1 vccd1 _11031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _11776_/CLK _10815_/D vssd1 vssd1 vccd1 vccd1 _10815_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11795_ _11801_/CLK _11795_/D vssd1 vssd1 vccd1 vccd1 _11795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10746_ _10765_/CLK _10746_/D vssd1 vssd1 vccd1 vccd1 _10746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ _10765_/CLK _10677_/D vssd1 vssd1 vccd1 vccd1 _10677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput208 _05483_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_4
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11229_ _11629_/CLK _11229_/D vssd1 vssd1 vccd1 vccd1 _11229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06770_ _11621_/Q _06704_/B _06769_/X vssd1 vssd1 vccd1 vccd1 _10243_/D sky130_fd_sc_hd__a21o_1
XFILLER_49_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05721_ _10974_/Q _05518_/Y _05524_/Y _10965_/Q vssd1 vssd1 vccd1 vccd1 _05721_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08440_ _11061_/Q _08436_/Y _08439_/Y _08440_/B2 vssd1 vssd1 vccd1 vccd1 _11061_/D
+ sky130_fd_sc_hd__a22o_1
X_05652_ _11287_/Q _05531_/Y _05555_/Y _11296_/Q _05651_/X vssd1 vssd1 vccd1 vccd1
+ _05652_/X sky130_fd_sc_hd__a221o_1
XFILLER_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05583_ _05619_/A1 _11388_/Q _11384_/Q _05619_/B2 _05581_/X vssd1 vssd1 vccd1 vccd1
+ _05583_/X sky130_fd_sc_hd__a221o_1
X_08371_ _10185_/A0 _08439_/B _08370_/X _08662_/C1 vssd1 vssd1 vccd1 vccd1 _11027_/D
+ sky130_fd_sc_hd__o211a_1
X_07322_ _08902_/B _08164_/B vssd1 vssd1 vccd1 vccd1 _07322_/Y sky130_fd_sc_hd__nor2_4
XFILLER_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07253_ _07254_/A _07854_/B vssd1 vssd1 vccd1 vccd1 _09175_/B sky130_fd_sc_hd__nor2_8
XFILLER_121_1320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06204_ _11319_/Q _06738_/A2 _06718_/C1 _06203_/X vssd1 vssd1 vccd1 vccd1 _06204_/X
+ sky130_fd_sc_hd__o211a_1
X_07184_ _10353_/Q _09228_/B vssd1 vssd1 vccd1 vccd1 _07184_/X sky130_fd_sc_hd__or2_1
XFILLER_145_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06135_ _11092_/Q _06629_/B1 _06133_/X _06134_/X vssd1 vssd1 vccd1 vccd1 _06135_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06066_ _10863_/Q _06455_/A2 _06412_/B1 _10836_/Q vssd1 vssd1 vccd1 vccd1 _06066_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout402 _05412_/Y vssd1 vssd1 vccd1 vccd1 _09571_/D sky130_fd_sc_hd__buf_6
XFILLER_87_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout413 _05357_/Y vssd1 vssd1 vccd1 vccd1 _09878_/B1 sky130_fd_sc_hd__buf_4
XFILLER_120_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout424 _05291_/Y vssd1 vssd1 vccd1 vccd1 _09565_/B sky130_fd_sc_hd__buf_8
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout435 _05238_/X vssd1 vssd1 vccd1 vccd1 _09875_/B1 sky130_fd_sc_hd__buf_4
XFILLER_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout446 _09909_/A2 vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout457 _05113_/Y vssd1 vssd1 vccd1 vccd1 _09876_/A2 sky130_fd_sc_hd__buf_4
X_09825_ _09825_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _11655_/D sky130_fd_sc_hd__and2_1
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout468 _07018_/B vssd1 vssd1 vccd1 vccd1 _09022_/C1 sky130_fd_sc_hd__buf_6
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout479 _07205_/A vssd1 vssd1 vccd1 vccd1 _07141_/B sky130_fd_sc_hd__buf_4
XFILLER_41_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09756_ _10551_/Q _09876_/A2 _09881_/B1 _10536_/Q _09755_/X vssd1 vssd1 vccd1 vccd1
+ _09757_/D sky130_fd_sc_hd__a221o_1
XFILLER_74_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06968_ _11608_/Q _09538_/C _06944_/A _09668_/C vssd1 vssd1 vccd1 vccd1 _06968_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08707_ _08947_/A1 _11208_/Q _08707_/S vssd1 vssd1 vccd1 vccd1 _08708_/B sky130_fd_sc_hd__mux2_1
X_05919_ _11315_/Q _08907_/A _08855_/A _11287_/Q _06718_/C1 vssd1 vssd1 vccd1 vccd1
+ _05922_/A sky130_fd_sc_hd__o221a_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09687_ _05393_/S _09682_/B _09682_/Y _11636_/Q _09686_/X vssd1 vssd1 vccd1 vccd1
+ _09688_/B sky130_fd_sc_hd__o221a_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ _10216_/Q _09447_/B vssd1 vssd1 vccd1 vccd1 _06899_/X sky130_fd_sc_hd__or2_4
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08638_ _08092_/X _08146_/S _08637_/X _08427_/A vssd1 vssd1 vccd1 vccd1 _11173_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _11139_/Q _07021_/A _08577_/S vssd1 vssd1 vccd1 vccd1 _08570_/B sky130_fd_sc_hd__mux2_1
X_10600_ _11781_/CLK _10600_/D vssd1 vssd1 vccd1 vccd1 _10600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11580_ _11584_/CLK _11580_/D vssd1 vssd1 vccd1 vccd1 _11580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10531_ _11745_/CLK _10531_/D vssd1 vssd1 vccd1 vccd1 _10531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10462_ _11136_/CLK _10462_/D vssd1 vssd1 vccd1 vccd1 _10462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10393_ _11720_/CLK _10393_/D vssd1 vssd1 vccd1 vccd1 _10393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11014_ _11756_/CLK _11014_/D vssd1 vssd1 vccd1 vccd1 _11014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout980 _10161_/A1 vssd1 vssd1 vccd1 vccd1 _09111_/A1 sky130_fd_sc_hd__buf_6
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout991 _07298_/B vssd1 vssd1 vccd1 vccd1 _11869_/A sky130_fd_sc_hd__clkbuf_16
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1082 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1082/HI io_oeb[12] sky130_fd_sc_hd__conb_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1093 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1093/HI io_oeb[23] sky130_fd_sc_hd__conb_1
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11778_ _11779_/CLK _11778_/D vssd1 vssd1 vccd1 vccd1 _11778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10729_ _11711_/CLK _10729_/D vssd1 vssd1 vccd1 vccd1 _10729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07940_ _10159_/A _08230_/B _10159_/C vssd1 vssd1 vccd1 vccd1 _08083_/S sky130_fd_sc_hd__or3_4
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11803_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07871_ _08789_/A1 _10754_/Q _07871_/S vssd1 vssd1 vccd1 vccd1 _07872_/B sky130_fd_sc_hd__mux2_1
XFILLER_151_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09610_ _10395_/Q _09567_/A _09570_/A _10627_/Q vssd1 vssd1 vccd1 vccd1 _09610_/X
+ sky130_fd_sc_hd__a22o_1
X_06822_ _10494_/Q _06872_/A2 _06818_/X _06821_/X vssd1 vssd1 vccd1 vccd1 _06822_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09541_ _09539_/X _09661_/B _09959_/B vssd1 vssd1 vccd1 vccd1 _09541_/Y sky130_fd_sc_hd__a21oi_4
X_06753_ _06744_/X _06747_/X _06752_/X vssd1 vssd1 vccd1 vccd1 _06753_/X sky130_fd_sc_hd__a21o_1
XFILLER_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05704_ _05704_/A _05704_/B _05704_/C vssd1 vssd1 vccd1 vccd1 _05704_/X sky130_fd_sc_hd__or3_4
XFILLER_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09472_ _09441_/B input25/X _09441_/A vssd1 vssd1 vccd1 vccd1 _09472_/X sky130_fd_sc_hd__o21a_1
X_06684_ _11616_/Q _06683_/X _06883_/B vssd1 vssd1 vccd1 vccd1 _10238_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08423_ _08423_/A1 _08383_/X _08422_/X _08947_/C1 vssd1 vssd1 vccd1 vccd1 _11052_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05635_ _11331_/Q _05591_/Y _05633_/Y _11314_/Q _05634_/X vssd1 vssd1 vccd1 vccd1
+ _05644_/A sky130_fd_sc_hd__a221o_1
XFILLER_24_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08354_ _08970_/A1 _11020_/Q _08354_/S vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__mux2_1
X_05566_ _11798_/Q _05076_/A _05079_/A _11792_/Q _05565_/X vssd1 vssd1 vccd1 vccd1
+ _05567_/B sky130_fd_sc_hd__a221o_4
XFILLER_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07305_ _08438_/A _08762_/B vssd1 vssd1 vccd1 vccd1 _07305_/Y sky130_fd_sc_hd__nor2_2
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05497_ _10242_/Q input54/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05497_/X sky130_fd_sc_hd__mux2_1
X_08285_ _08423_/A1 _08276_/S _08284_/X _08921_/C1 vssd1 vssd1 vccd1 vccd1 _10974_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07236_ _07235_/X _10386_/Q _07246_/S vssd1 vssd1 vccd1 vccd1 _10386_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07167_ _09129_/A1 _07172_/S _07166_/X _07884_/C1 vssd1 vssd1 vccd1 vccd1 _10344_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06118_ _11108_/Q _06716_/A2 _06716_/B1 _11244_/Q vssd1 vssd1 vccd1 vccd1 _06119_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07098_ _07617_/A _07098_/B vssd1 vssd1 vccd1 vccd1 _07098_/X sky130_fd_sc_hd__or2_1
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06049_ _06040_/X _06042_/X _06043_/X _06048_/X vssd1 vssd1 vccd1 vccd1 _06049_/X
+ sky130_fd_sc_hd__a31o_2
Xfanout221 _07338_/Y vssd1 vssd1 vccd1 vccd1 _07346_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout232 _07491_/S vssd1 vssd1 vccd1 vccd1 _07496_/S sky130_fd_sc_hd__buf_6
XFILLER_119_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout243 _09488_/Y vssd1 vssd1 vccd1 vccd1 _09500_/B sky130_fd_sc_hd__buf_2
XFILLER_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout254 _08683_/S vssd1 vssd1 vccd1 vccd1 _08707_/S sky130_fd_sc_hd__buf_8
Xfanout265 _08383_/X vssd1 vssd1 vccd1 vccd1 _08404_/S sky130_fd_sc_hd__clkbuf_16
Xfanout276 _08097_/X vssd1 vssd1 vccd1 vccd1 _08360_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout287 _07893_/B vssd1 vssd1 vccd1 vccd1 _07901_/B sky130_fd_sc_hd__buf_4
X_09808_ _10524_/Q _09568_/B _09568_/C _10526_/Q _09802_/X vssd1 vssd1 vccd1 vccd1
+ _09811_/B sky130_fd_sc_hd__a221o_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout298 _07638_/X vssd1 vssd1 vccd1 vccd1 _08102_/S sky130_fd_sc_hd__buf_6
Xclkbuf_4_15__f_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_77_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09739_ _09739_/A _09739_/B _09739_/C _09739_/D vssd1 vssd1 vccd1 vccd1 _09740_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11701_ _11744_/CLK _11701_/D vssd1 vssd1 vccd1 vccd1 _11701_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11632_/CLK _11632_/D vssd1 vssd1 vccd1 vccd1 _11632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11563_ _11810_/CLK _11563_/D vssd1 vssd1 vccd1 vccd1 _11563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10514_ _10725_/CLK _10514_/D vssd1 vssd1 vccd1 vccd1 _10514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11494_ _11497_/CLK _11494_/D vssd1 vssd1 vccd1 vccd1 _11494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ _11780_/CLK _10445_/D vssd1 vssd1 vccd1 vccd1 _10445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10376_ _11744_/CLK _10376_/D vssd1 vssd1 vccd1 vccd1 _10376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 _05692_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _10086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_192 _07059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05420_ _11238_/Q _11237_/Q _05471_/A vssd1 vssd1 vccd1 vccd1 _05422_/C sky130_fd_sc_hd__mux2_1
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05351_ _11310_/Q _11309_/Q _05385_/S vssd1 vssd1 vccd1 vccd1 _05356_/C sky130_fd_sc_hd__mux2_1
XFILLER_81_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05282_ _10896_/Q _10895_/Q _05430_/S vssd1 vssd1 vccd1 vccd1 _05282_/X sky130_fd_sc_hd__mux2_1
X_08070_ _08469_/A _08427_/B _08069_/X _08351_/C1 vssd1 vssd1 vccd1 vccd1 _10860_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07021_ _07021_/A _07107_/B vssd1 vssd1 vccd1 vccd1 _07022_/B sky130_fd_sc_hd__and2_4
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08972_ _08972_/A _09271_/B _09038_/C vssd1 vssd1 vccd1 vccd1 _08972_/X sky130_fd_sc_hd__or3_4
XFILLER_102_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07923_ _08939_/A1 _10779_/Q _09218_/S vssd1 vssd1 vccd1 vccd1 _07924_/B sky130_fd_sc_hd__mux2_1
XFILLER_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07854_ _07854_/A _07854_/B vssd1 vssd1 vccd1 vccd1 _07854_/X sky130_fd_sc_hd__or2_1
XFILLER_69_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06805_ _11472_/Q _07152_/A _06805_/B1 _10551_/Q vssd1 vssd1 vccd1 vccd1 _06805_/X
+ sky130_fd_sc_hd__o22a_1
X_07785_ _07785_/A0 _10700_/Q _07817_/S vssd1 vssd1 vccd1 vccd1 _07786_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09524_ _09502_/A _09489_/C _09495_/C _11618_/Q vssd1 vssd1 vccd1 vccd1 _09526_/B
+ sky130_fd_sc_hd__a31o_1
X_06736_ _11208_/Q _06736_/A2 _08765_/A _11258_/Q vssd1 vssd1 vccd1 vccd1 _06736_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09441_/B input12/X _09441_/Y input29/X _09454_/X vssd1 vssd1 vccd1 vccd1
+ _09455_/X sky130_fd_sc_hd__a221o_1
X_06667_ _10388_/Q _06860_/A2 _07539_/A _10325_/Q _06666_/X vssd1 vssd1 vccd1 vccd1
+ _06667_/X sky130_fd_sc_hd__o221a_1
X_08406_ _08789_/A1 _11044_/Q _08414_/S vssd1 vssd1 vccd1 vccd1 _08407_/B sky130_fd_sc_hd__mux2_1
X_05618_ _05618_/A1 _11372_/Q _11369_/Q _11624_/Q _05616_/X vssd1 vssd1 vccd1 vccd1
+ _05621_/A sky130_fd_sc_hd__a221o_4
X_09386_ _10114_/A0 _11553_/Q _09390_/S vssd1 vssd1 vccd1 vccd1 _11553_/D sky130_fd_sc_hd__mux2_1
X_06598_ _10886_/Q _06468_/B _06152_/B _10933_/Q _06597_/X vssd1 vssd1 vccd1 vccd1
+ _06598_/X sky130_fd_sc_hd__o221a_1
XFILLER_61_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08337_ _09999_/A0 _08360_/S _08336_/X _08351_/C1 vssd1 vssd1 vccd1 vccd1 _11011_/D
+ sky130_fd_sc_hd__o211a_1
X_05549_ _05549_/A _05549_/B vssd1 vssd1 vccd1 vccd1 _05549_/Y sky130_fd_sc_hd__nor2_8
XFILLER_138_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08268_ _08789_/A1 _10966_/Q _08272_/S vssd1 vssd1 vccd1 vccd1 _08269_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ _07147_/A _07204_/B _07771_/B1 _10376_/Q vssd1 vssd1 vccd1 vccd1 _10376_/D
+ sky130_fd_sc_hd__a22o_1
X_08199_ _10158_/A _08649_/C _09037_/C vssd1 vssd1 vccd1 vccd1 _08902_/C sky130_fd_sc_hd__and3_4
X_10230_ _11628_/CLK _10230_/D vssd1 vssd1 vccd1 vccd1 _10230_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10161_ _10161_/A1 _10159_/X _10160_/X _10175_/C1 vssd1 vssd1 vccd1 vccd1 _11792_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1005 input79/X vssd1 vssd1 vccd1 vccd1 _05745_/A sky130_fd_sc_hd__buf_8
Xfanout1016 _10105_/A1 vssd1 vssd1 vccd1 vccd1 _10117_/A0 sky130_fd_sc_hd__buf_2
Xfanout1027 _10175_/A1 vssd1 vssd1 vccd1 vccd1 _08987_/A1 sky130_fd_sc_hd__buf_6
XFILLER_134_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10092_ _10142_/A1 _10104_/B _10156_/B1 vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__a21o_1
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1038 _09971_/A0 vssd1 vssd1 vccd1 vccd1 _10114_/A0 sky130_fd_sc_hd__buf_4
XFILLER_43_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1049 input112/X vssd1 vssd1 vccd1 vccd1 _07092_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_75_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10994_ _11756_/CLK _10994_/D vssd1 vssd1 vccd1 vccd1 _10994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11615_ _11663_/CLK _11615_/D vssd1 vssd1 vccd1 vccd1 _11615_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_156_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11546_ _11800_/CLK _11546_/D vssd1 vssd1 vccd1 vccd1 _11546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11477_ _11477_/CLK _11477_/D vssd1 vssd1 vccd1 vccd1 _11477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10428_ _11628_/CLK _10428_/D vssd1 vssd1 vccd1 vccd1 _10428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10359_ _11710_/CLK _10359_/D vssd1 vssd1 vccd1 vccd1 _10359_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07570_ _10056_/A _07570_/B vssd1 vssd1 vccd1 vccd1 _10568_/D sky130_fd_sc_hd__or2_1
XFILLER_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06521_ _10346_/Q _06649_/A2 _06517_/X _06520_/X vssd1 vssd1 vccd1 vccd1 _06521_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09240_ input104/X _11472_/Q _09240_/S vssd1 vssd1 vccd1 vccd1 _09240_/X sky130_fd_sc_hd__mux2_1
X_06452_ _11610_/Q _06665_/A2 _06450_/X _06622_/B2 _06451_/X vssd1 vssd1 vccd1 vccd1
+ _10232_/D sky130_fd_sc_hd__a221o_1
XFILLER_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05403_ _10586_/Q _10585_/Q _09538_/A vssd1 vssd1 vccd1 vccd1 _05406_/B sky130_fd_sc_hd__mux2_1
X_09171_ _11430_/Q _09171_/B vssd1 vssd1 vccd1 vccd1 _09171_/X sky130_fd_sc_hd__or2_1
X_06383_ _11064_/Q _06629_/A2 _06453_/B1 _10642_/Q vssd1 vssd1 vccd1 vccd1 _06387_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08122_ _09976_/A _08649_/C _09037_/C vssd1 vssd1 vccd1 vccd1 _08637_/C sky130_fd_sc_hd__and3_4
X_05334_ _05334_/A _05334_/B _05334_/C _05334_/D vssd1 vssd1 vccd1 vccd1 _05335_/B
+ sky130_fd_sc_hd__or4_4
X_08053_ _09358_/A _08649_/C _09037_/C vssd1 vssd1 vccd1 vccd1 _08426_/B sky130_fd_sc_hd__and3_4
XFILLER_107_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05265_ _10436_/Q _10435_/Q _05391_/S vssd1 vssd1 vccd1 vccd1 _05269_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07004_ _09668_/A _08847_/A vssd1 vssd1 vccd1 vccd1 _07004_/Y sky130_fd_sc_hd__nand2_4
XFILLER_66_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05196_ _11030_/Q _11029_/Q _05414_/S vssd1 vssd1 vccd1 vccd1 _05196_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput108 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 _07039_/A sky130_fd_sc_hd__buf_4
X_08955_ _08955_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _09491_/C sky130_fd_sc_hd__or2_1
XFILLER_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput119 wbs_we_i vssd1 vssd1 vccd1 vccd1 _05819_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07906_ _07916_/A _07906_/B vssd1 vssd1 vccd1 vccd1 _10770_/D sky130_fd_sc_hd__or2_1
XFILLER_102_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08886_ _08939_/A1 _11300_/Q _08890_/S vssd1 vssd1 vccd1 vccd1 _08887_/B sky130_fd_sc_hd__mux2_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07837_ _07034_/A _07820_/B _07821_/A _10732_/Q vssd1 vssd1 vccd1 vccd1 _10732_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07768_ _10688_/Q _07232_/X _07773_/S vssd1 vssd1 vccd1 vccd1 _10688_/D sky130_fd_sc_hd__mux2_1
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09507_ _09515_/B _09515_/C _09511_/C vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__and3b_1
XFILLER_53_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06719_ _11207_/Q _06719_/A2 _09038_/A _11170_/Q _06718_/X vssd1 vssd1 vccd1 vccd1
+ _06720_/B sky130_fd_sc_hd__o221a_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ _10647_/Q _07694_/Y _07696_/Y _07309_/X vssd1 vssd1 vccd1 vccd1 _10647_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _11591_/Q _11650_/Q _09440_/S vssd1 vssd1 vccd1 vccd1 _11591_/D sky130_fd_sc_hd__mux2_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _10168_/A1 _09359_/X _09368_/X _09995_/C1 vssd1 vssd1 vccd1 vccd1 _11542_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11400_ _11462_/CLK _11400_/D vssd1 vssd1 vccd1 vccd1 _11400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_70 _05668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_81 _11587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11331_ _11393_/CLK _11331_/D vssd1 vssd1 vccd1 vccd1 _11331_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_92 _09950_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11262_ _11262_/CLK _11262_/D vssd1 vssd1 vccd1 vccd1 _11262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10213_ _11634_/CLK _10213_/D vssd1 vssd1 vccd1 vccd1 _10213_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11193_ _11251_/CLK _11193_/D vssd1 vssd1 vccd1 vccd1 _11193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10144_ _11785_/Q _10154_/B vssd1 vssd1 vccd1 vccd1 _10144_/X sky130_fd_sc_hd__or2_1
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10075_ _10111_/A0 _11735_/Q _10082_/S vssd1 vssd1 vccd1 vccd1 _11735_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ _11136_/CLK _10977_/D vssd1 vssd1 vccd1 vccd1 _10977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11529_ _11735_/CLK _11529_/D vssd1 vssd1 vccd1 vccd1 _11529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout809 _06766_/A2 vssd1 vssd1 vccd1 vccd1 _07153_/A sky130_fd_sc_hd__buf_6
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08740_ _11227_/Q _08750_/B vssd1 vssd1 vccd1 vccd1 _08740_/X sky130_fd_sc_hd__or2_1
XFILLER_100_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05952_ _11521_/Q _09326_/A _08245_/A _11481_/Q vssd1 vssd1 vccd1 vccd1 _05952_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08671_ _09114_/A1 _11190_/Q _08707_/S vssd1 vssd1 vccd1 vccd1 _08672_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05883_ _07082_/A _05881_/X _05882_/X _05816_/A vssd1 vssd1 vccd1 vccd1 _05883_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_94_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07622_ _10596_/Q _07613_/A _08037_/B _07621_/X vssd1 vssd1 vccd1 vccd1 _10596_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07553_ _10021_/A0 _10560_/Q _07593_/S vssd1 vssd1 vccd1 vccd1 _07554_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06504_ _11235_/Q _06541_/A2 _06504_/B1 _11009_/Q _06503_/X vssd1 vssd1 vccd1 vccd1
+ _06504_/X sky130_fd_sc_hd__o221a_1
X_07484_ _10026_/A _07484_/B vssd1 vssd1 vccd1 vccd1 _10520_/D sky130_fd_sc_hd__or2_1
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09223_ _11461_/Q _09205_/Y _09209_/Y _07451_/X vssd1 vssd1 vccd1 vccd1 _11461_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06435_ _10539_/Q _09109_/A _06434_/X _06873_/D1 vssd1 vssd1 vccd1 vccd1 _06435_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09154_ _09154_/A _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09154_/X sky130_fd_sc_hd__or3_4
X_06366_ _10402_/Q _06804_/B _06806_/A2 _10563_/Q vssd1 vssd1 vccd1 vccd1 _06366_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08105_ _10877_/Q _08120_/S _07642_/S _07229_/B vssd1 vssd1 vccd1 vccd1 _10877_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05317_ _10878_/Q _10877_/Q _05393_/S vssd1 vssd1 vccd1 vccd1 _05318_/D sky130_fd_sc_hd__mux2_1
X_09085_ _09275_/A1 _09099_/B _08873_/A vssd1 vssd1 vccd1 vccd1 _09085_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06297_ _11546_/Q _09359_/A _09977_/A _11684_/Q _06297_/C1 vssd1 vssd1 vccd1 vccd1
+ _06297_/X sky130_fd_sc_hd__o221a_1
XFILLER_120_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08036_ _08851_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _10842_/D sky130_fd_sc_hd__or2_1
Xinput90 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__buf_8
X_05248_ _05248_/A _05248_/B _05248_/C _05248_/D vssd1 vssd1 vccd1 vccd1 _05248_/Y
+ sky130_fd_sc_hd__nor4_4
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05179_ _05179_/A _05179_/B vssd1 vssd1 vccd1 vccd1 _05179_/Y sky130_fd_sc_hd__nor2_8
XFILLER_107_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09987_ _10168_/A1 _09977_/X _09986_/X _09993_/C1 vssd1 vssd1 vccd1 vccd1 _11680_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08938_ _11328_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08938_/X sky130_fd_sc_hd__or2_1
XFILLER_130_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08869_ _08869_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _11291_/D sky130_fd_sc_hd__or2_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ _11601_/CLK _10900_/D vssd1 vssd1 vccd1 vccd1 _10900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10831_ _11604_/CLK _10831_/D vssd1 vssd1 vccd1 vccd1 _10831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10762_ _10782_/CLK _10762_/D vssd1 vssd1 vccd1 vccd1 _10762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10693_ _10725_/CLK _10693_/D vssd1 vssd1 vccd1 vccd1 _10693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ _11393_/CLK _11314_/D vssd1 vssd1 vccd1 vccd1 _11314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11245_ _11319_/CLK _11245_/D vssd1 vssd1 vccd1 vccd1 _11245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11176_ _11177_/CLK _11176_/D vssd1 vssd1 vccd1 vccd1 _11176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10127_ _07018_/A _11773_/Q _10135_/S vssd1 vssd1 vccd1 vccd1 _11773_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10058_ _10058_/A _10058_/B vssd1 vssd1 vccd1 vccd1 _11720_/D sky130_fd_sc_hd__or2_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_69_wb_clk_i clkbuf_leaf_69_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11428_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06220_ _11495_/Q _06738_/A2 _06717_/B1 _11346_/Q vssd1 vssd1 vccd1 vccd1 _06220_/X
+ sky130_fd_sc_hd__o22a_1
X_06151_ _06151_/A _06151_/B _06151_/C vssd1 vssd1 vccd1 vccd1 _06151_/X sky130_fd_sc_hd__and3_1
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05102_ _05729_/A input87/X vssd1 vssd1 vccd1 vccd1 _10255_/D sky130_fd_sc_hd__and2_4
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06082_ _06663_/A _10227_/Q vssd1 vssd1 vccd1 vccd1 _06082_/X sky130_fd_sc_hd__and2_1
XFILLER_145_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09910_ _10493_/Q _09571_/A _09567_/A _10495_/Q _09909_/X vssd1 vssd1 vccd1 vccd1
+ _09917_/A sky130_fd_sc_hd__a221o_1
XFILLER_125_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout606 _06430_/A2 vssd1 vssd1 vccd1 vccd1 _06308_/A2 sky130_fd_sc_hd__buf_4
Xfanout617 _06748_/A2 vssd1 vssd1 vccd1 vccd1 _06106_/B sky130_fd_sc_hd__buf_2
X_09841_ _11454_/Q _09873_/A2 _09571_/D _10771_/Q _09840_/X vssd1 vssd1 vccd1 vccd1
+ _09842_/D sky130_fd_sc_hd__a221o_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout628 _05736_/Y vssd1 vssd1 vccd1 vccd1 _09325_/A sky130_fd_sc_hd__buf_12
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout639 _05079_/Y vssd1 vssd1 vccd1 vccd1 _05620_/B2 sky130_fd_sc_hd__clkbuf_16
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _05427_/S _09672_/B _09674_/A _11588_/Q vssd1 vssd1 vccd1 vccd1 _09772_/X
+ sky130_fd_sc_hd__o22a_1
X_06984_ _09256_/A1 _06976_/X _06983_/X _06990_/C1 vssd1 vssd1 vccd1 vccd1 _10259_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _11218_/Q _08726_/S _07852_/S _08817_/B2 vssd1 vssd1 vccd1 vccd1 _11218_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05935_ _11233_/Q _06541_/A2 _06504_/B1 _11002_/Q vssd1 vssd1 vccd1 vccd1 _05935_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08654_ _07005_/A _08750_/B _08653_/X vssd1 vssd1 vccd1 vccd1 _11182_/D sky130_fd_sc_hd__a21o_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05866_ _10910_/Q _08166_/A _06513_/A2 _10436_/Q _05865_/X vssd1 vssd1 vccd1 vccd1
+ _05866_/X sky130_fd_sc_hd__o221a_1
XFILLER_96_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07605_ _10585_/Q _07597_/Y _07600_/Y _07016_/X vssd1 vssd1 vccd1 vccd1 _10585_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _07104_/A _11148_/Q _08589_/S vssd1 vssd1 vccd1 vccd1 _08586_/B sky130_fd_sc_hd__mux2_1
X_05797_ _11123_/Q _07222_/A _05796_/X _06550_/C1 vssd1 vssd1 vccd1 vccd1 _05797_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07536_ _07934_/A _07536_/B vssd1 vssd1 vccd1 vccd1 _10552_/D sky130_fd_sc_hd__or2_1
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07467_ _07059_/A _10511_/Q _07477_/S vssd1 vssd1 vccd1 vccd1 _07468_/B sky130_fd_sc_hd__mux2_1
X_09206_ _09206_/A _09206_/B vssd1 vssd1 vccd1 vccd1 _09206_/Y sky130_fd_sc_hd__nand2_2
XFILLER_139_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06418_ _10855_/Q _08054_/A _06416_/X _06417_/X vssd1 vssd1 vccd1 vccd1 _06418_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07398_ _07476_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _10475_/D sky130_fd_sc_hd__or2_1
XFILLER_124_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09137_ _09276_/A1 _09149_/B _09173_/B1 vssd1 vssd1 vccd1 vccd1 _09137_/X sky130_fd_sc_hd__a21o_1
X_06349_ _11368_/Q _09016_/A _08994_/A _11358_/Q _06349_/C1 vssd1 vssd1 vccd1 vccd1
+ _06349_/X sky130_fd_sc_hd__o221a_1
XFILLER_120_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09068_ _11382_/Q _09060_/X _09067_/X vssd1 vssd1 vccd1 vccd1 _11382_/D sky130_fd_sc_hd__a21o_1
XFILLER_118_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08019_ _10834_/Q _08037_/B vssd1 vssd1 vccd1 vccd1 _08019_/X sky130_fd_sc_hd__or2_1
XFILLER_104_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11030_ _11067_/CLK _11030_/D vssd1 vssd1 vccd1 vccd1 _11030_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _11776_/CLK _10814_/D vssd1 vssd1 vccd1 vccd1 _10814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _11800_/CLK _11794_/D vssd1 vssd1 vccd1 vccd1 _11794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ _11770_/CLK _10745_/D vssd1 vssd1 vccd1 vccd1 _10745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10676_ _10785_/CLK _10676_/D vssd1 vssd1 vccd1 vccd1 _10676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput209 _05484_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_4
XFILLER_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_116_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11720_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11228_ _11629_/CLK _11228_/D vssd1 vssd1 vccd1 vccd1 _11228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11159_ _11329_/CLK _11159_/D vssd1 vssd1 vccd1 vccd1 _11159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05720_ _10970_/Q _05561_/Y _05585_/Y _10969_/Q _05719_/X vssd1 vssd1 vccd1 vccd1
+ _05728_/A sky130_fd_sc_hd__a221o_1
XFILLER_82_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05651_ _11288_/Q _05567_/Y _05621_/Y _11297_/Q vssd1 vssd1 vccd1 vccd1 _05651_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _11027_/Q _08438_/B vssd1 vssd1 vccd1 vccd1 _08370_/X sky130_fd_sc_hd__or2_1
X_05582_ _05618_/A1 _11382_/Q _11379_/Q _05606_/B2 _05580_/X vssd1 vssd1 vccd1 vccd1
+ _05585_/A sky130_fd_sc_hd__a221o_4
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07321_ _09293_/A _08665_/C _10159_/C vssd1 vssd1 vccd1 vccd1 _08162_/S sky130_fd_sc_hd__or3_4
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07252_ _10395_/Q _07249_/S _07251_/X _09206_/A vssd1 vssd1 vccd1 vccd1 _10395_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06203_ _11039_/Q _06735_/A2 _06739_/A2 _11291_/Q _06202_/X vssd1 vssd1 vccd1 vccd1
+ _06203_/X sky130_fd_sc_hd__o221a_1
XFILLER_121_1332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07183_ _10043_/A _07183_/B vssd1 vssd1 vccd1 vccd1 _10352_/D sky130_fd_sc_hd__or2_1
XFILLER_30_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06134_ _11058_/Q _08054_/A _06632_/A2 _10892_/Q _06392_/C1 vssd1 vssd1 vccd1 vccd1
+ _06134_/X sky130_fd_sc_hd__o221a_1
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06065_ _10419_/Q _06318_/A2 _06589_/A2 _11003_/Q vssd1 vssd1 vccd1 vccd1 _06065_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout403 _05412_/Y vssd1 vssd1 vccd1 vccd1 _09872_/B1 sky130_fd_sc_hd__buf_4
XFILLER_154_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout414 _05346_/Y vssd1 vssd1 vccd1 vccd1 _09950_/B1 sky130_fd_sc_hd__buf_8
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout425 _05291_/Y vssd1 vssd1 vccd1 vccd1 _09884_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout436 _05224_/Y vssd1 vssd1 vccd1 vccd1 _09568_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout447 _05168_/Y vssd1 vssd1 vccd1 vccd1 _09909_/A2 sky130_fd_sc_hd__buf_6
X_09824_ _09522_/B _09823_/Y _09824_/S vssd1 vssd1 vccd1 vccd1 _09825_/B sky130_fd_sc_hd__mux2_1
XFILLER_154_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout458 _06938_/B vssd1 vssd1 vccd1 vccd1 _09681_/B sky130_fd_sc_hd__buf_6
XFILLER_28_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout469 _08662_/C1 vssd1 vssd1 vccd1 vccd1 _08753_/C1 sky130_fd_sc_hd__buf_6
XFILLER_101_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_14__f_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_85_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09755_ _10545_/Q _09881_/A2 _09565_/C _10543_/Q vssd1 vssd1 vccd1 vccd1 _09755_/X
+ sky130_fd_sc_hd__a22o_1
X_06967_ _06967_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09668_/C sky130_fd_sc_hd__nand2_4
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05918_ _05912_/X _05917_/X _07151_/B vssd1 vssd1 vccd1 vccd1 _05918_/X sky130_fd_sc_hd__o21a_2
X_08706_ _08893_/A1 _08707_/S _08705_/X _09078_/C1 vssd1 vssd1 vccd1 vccd1 _11207_/D
+ sky130_fd_sc_hd__o211a_1
X_09686_ _11640_/Q _09692_/B vssd1 vssd1 vccd1 vccd1 _09686_/X sky130_fd_sc_hd__or2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06898_ _10216_/Q _09447_/B vssd1 vssd1 vccd1 vccd1 _06898_/Y sky130_fd_sc_hd__nor2_8
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _11173_/Q _08902_/B _08637_/C vssd1 vssd1 vccd1 vccd1 _08637_/X sky130_fd_sc_hd__or3_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05849_ _10655_/Q _07455_/A vssd1 vssd1 vccd1 vccd1 _05849_/X sky130_fd_sc_hd__or2_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _08733_/A _08568_/B vssd1 vssd1 vccd1 vccd1 _11138_/D sky130_fd_sc_hd__or2_1
XFILLER_23_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07519_ _07211_/A _10544_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _07520_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08499_ _11100_/Q _08503_/B vssd1 vssd1 vccd1 vccd1 _08499_/X sky130_fd_sc_hd__or2_1
X_10530_ _10735_/CLK _10530_/D vssd1 vssd1 vccd1 vccd1 _10530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10461_ _11308_/CLK _10461_/D vssd1 vssd1 vccd1 vccd1 _10461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10392_ _11706_/CLK _10392_/D vssd1 vssd1 vccd1 vccd1 _10392_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11013_ _11756_/CLK _11013_/D vssd1 vssd1 vccd1 vccd1 _11013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout970 _08931_/A1 vssd1 vssd1 vccd1 vccd1 _08789_/A1 sky130_fd_sc_hd__buf_6
XFILLER_93_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout981 _07303_/A vssd1 vssd1 vccd1 vccd1 _10161_/A1 sky130_fd_sc_hd__buf_8
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout992 _07690_/B vssd1 vssd1 vccd1 vccd1 _06344_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapped_tms1x00_1083 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1083/HI io_oeb[13] sky130_fd_sc_hd__conb_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1094 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1094/HI io_oeb[24] sky130_fd_sc_hd__conb_1
XFILLER_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11777_ _11777_/CLK _11777_/D vssd1 vssd1 vccd1 vccd1 _11777_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10728_ _11743_/CLK _10728_/D vssd1 vssd1 vccd1 vccd1 _10728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ _10765_/CLK _10659_/D vssd1 vssd1 vccd1 vccd1 _10659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07870_ _09129_/A1 _07970_/S _07869_/X _07894_/C1 vssd1 vssd1 vccd1 vccd1 _10753_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06821_ _10394_/Q _06860_/A2 _06820_/X _06849_/C1 vssd1 vssd1 vccd1 vccd1 _06821_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09540_ _09540_/A _09668_/B _09668_/C _09668_/D vssd1 vssd1 vccd1 vccd1 _09661_/B
+ sky130_fd_sc_hd__or4_4
Xclkbuf_leaf_84_wb_clk_i clkbuf_leaf_85_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11329_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_06752_ _10411_/Q _07254_/A _06748_/X _06751_/X vssd1 vssd1 vccd1 vccd1 _06752_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_114_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11310_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_97_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05703_ _05703_/A _05703_/B _05703_/C vssd1 vssd1 vccd1 vccd1 _05704_/C sky130_fd_sc_hd__or3_1
X_09471_ _09680_/C _09475_/A _09470_/Y _09478_/A vssd1 vssd1 vccd1 vccd1 _11600_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06683_ _06852_/A3 _06676_/X _06681_/X _06682_/X vssd1 vssd1 vccd1 vccd1 _06683_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_110_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08422_ _11052_/Q _08422_/B vssd1 vssd1 vccd1 vccd1 _08422_/X sky130_fd_sc_hd__or2_1
X_05634_ _11318_/Q _05609_/Y _05627_/Y _11313_/Q vssd1 vssd1 vccd1 vccd1 _05634_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08353_ _08969_/A1 _08354_/S _08352_/X _08831_/C1 vssd1 vssd1 vccd1 vccd1 _11019_/D
+ sky130_fd_sc_hd__o211a_1
X_05565_ _11801_/Q _05619_/A1 _05619_/B2 _11797_/Q _05563_/X vssd1 vssd1 vccd1 vccd1
+ _05565_/X sky130_fd_sc_hd__a221o_1
XFILLER_20_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07304_ _10417_/Q _07302_/Y _07303_/X _08760_/S _08439_/A vssd1 vssd1 vccd1 vccd1
+ _10417_/D sky130_fd_sc_hd__o221a_1
X_08284_ _10974_/Q _08284_/B vssd1 vssd1 vccd1 vccd1 _08284_/X sky130_fd_sc_hd__or2_1
X_05496_ _10241_/Q input52/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05496_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07235_ _10134_/A0 _10028_/A _07333_/A vssd1 vssd1 vccd1 vccd1 _07235_/X sky130_fd_sc_hd__a21o_2
XFILLER_20_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07166_ _10344_/Q _09228_/B vssd1 vssd1 vccd1 vccd1 _07166_/X sky130_fd_sc_hd__or2_1
XFILLER_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06117_ _11038_/Q _06735_/A2 _06717_/B1 _10960_/Q vssd1 vssd1 vccd1 vccd1 _06119_/B
+ sky130_fd_sc_hd__o22a_1
X_07097_ _07022_/B _08645_/S _07086_/Y _10304_/Q _07318_/A vssd1 vssd1 vccd1 vccd1
+ _10304_/D sky130_fd_sc_hd__a221o_1
XFILLER_117_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06048_ _11454_/Q _06862_/A2 _06044_/X _06047_/X vssd1 vssd1 vccd1 vccd1 _06048_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout222 _07233_/S vssd1 vssd1 vccd1 vccd1 _07246_/S sky130_fd_sc_hd__buf_6
Xfanout233 _07047_/Y vssd1 vssd1 vccd1 vccd1 _07491_/S sky130_fd_sc_hd__buf_6
Xfanout244 _08945_/A2 vssd1 vssd1 vccd1 vccd1 _08940_/S sky130_fd_sc_hd__buf_4
Xfanout255 _08650_/X vssd1 vssd1 vccd1 vccd1 _08748_/S sky130_fd_sc_hd__buf_6
XFILLER_8_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout266 _08365_/X vssd1 vssd1 vccd1 vccd1 _08439_/B sky130_fd_sc_hd__buf_6
X_09807_ _10298_/Q _09567_/A _09571_/C _10528_/Q _09803_/X vssd1 vssd1 vccd1 vccd1
+ _09811_/A sky130_fd_sc_hd__a221o_1
XFILLER_8_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout277 _08097_/X vssd1 vssd1 vccd1 vccd1 _08354_/S sky130_fd_sc_hd__clkbuf_4
Xfanout288 _07893_/B vssd1 vssd1 vccd1 vccd1 _07883_/B sky130_fd_sc_hd__buf_4
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout299 _07630_/B vssd1 vssd1 vccd1 vccd1 _08820_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_28_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07999_ _09396_/A0 _10824_/Q _08015_/S vssd1 vssd1 vccd1 vccd1 _08000_/B sky130_fd_sc_hd__mux2_1
XFILLER_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09738_ _10345_/Q _09876_/B1 _09567_/C _10344_/Q _09737_/X vssd1 vssd1 vccd1 vccd1
+ _09739_/D sky130_fd_sc_hd__a221o_2
XFILLER_41_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _09959_/B _09669_/B vssd1 vssd1 vccd1 vccd1 _09669_/Y sky130_fd_sc_hd__nor2_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11703_/CLK _11700_/D vssd1 vssd1 vccd1 vccd1 _11700_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11702_/CLK _11631_/D vssd1 vssd1 vccd1 vccd1 _11631_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11562_ _11675_/CLK _11562_/D vssd1 vssd1 vccd1 vccd1 _11562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10513_ _11743_/CLK _10513_/D vssd1 vssd1 vccd1 vccd1 _10513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11493_ _11497_/CLK _11493_/D vssd1 vssd1 vccd1 vccd1 _11493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10444_ _11766_/CLK _10444_/D vssd1 vssd1 vccd1 vccd1 _10444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10375_ _11722_/CLK _10375_/D vssd1 vssd1 vccd1 vccd1 _10375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _10119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_182 _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_193 _08929_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05350_ _11144_/Q _11143_/Q _09680_/B vssd1 vssd1 vccd1 vccd1 _05356_/B sky130_fd_sc_hd__mux2_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_131_wb_clk_i clkbuf_4_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10727_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_05281_ _05281_/A _05281_/B vssd1 vssd1 vccd1 vccd1 _05281_/Y sky130_fd_sc_hd__nor2_8
XFILLER_88_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07020_ _10270_/Q _07019_/X _07038_/S vssd1 vssd1 vccd1 vccd1 _10270_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _08971_/A _10136_/B _09037_/C vssd1 vssd1 vccd1 vccd1 _08989_/B sky130_fd_sc_hd__and3_4
X_07922_ _07922_/A _07922_/B vssd1 vssd1 vccd1 vccd1 _10778_/D sky130_fd_sc_hd__or2_1
XFILLER_96_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07853_ _07853_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07853_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06804_ _11438_/Q _06804_/B vssd1 vssd1 vccd1 vccd1 _06804_/X sky130_fd_sc_hd__or2_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07784_ _08684_/A _07784_/B vssd1 vssd1 vccd1 vccd1 _10699_/D sky130_fd_sc_hd__or2_1
XFILLER_65_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09523_ _09825_/A _09523_/B _09523_/C vssd1 vssd1 vccd1 vccd1 _11617_/D sky130_fd_sc_hd__and3_1
X_06735_ _11052_/Q _06735_/A2 _06735_/B1 _11171_/Q vssd1 vssd1 vccd1 vccd1 _06735_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09454_ _09441_/B input20/X _09441_/A vssd1 vssd1 vccd1 vccd1 _09454_/X sky130_fd_sc_hd__o21a_1
X_06666_ _10273_/Q _06999_/A vssd1 vssd1 vccd1 vccd1 _06666_/X sky130_fd_sc_hd__or2_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05617_ _09552_/A1 _11377_/Q _11371_/Q _05078_/A vssd1 vssd1 vccd1 vccd1 _05617_/X
+ sky130_fd_sc_hd__a22o_1
X_08405_ _08781_/A _08405_/B vssd1 vssd1 vccd1 vccd1 _11043_/D sky130_fd_sc_hd__or2_1
X_09385_ _10113_/A0 _11552_/Q _09390_/S vssd1 vssd1 vccd1 vccd1 _11552_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06597_ _11231_/Q _08650_/A _06640_/B1 _11143_/Q vssd1 vssd1 vccd1 vccd1 _06597_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_75_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08336_ _11011_/Q _08362_/B vssd1 vssd1 vccd1 vccd1 _08336_/X sky130_fd_sc_hd__or2_1
X_05548_ _05076_/A _11494_/Q _11489_/Q _05620_/B2 _05547_/X vssd1 vssd1 vccd1 vccd1
+ _05549_/B sky130_fd_sc_hd__a221o_4
XFILLER_71_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08267_ _08781_/A _08267_/B vssd1 vssd1 vccd1 vccd1 _10965_/D sky130_fd_sc_hd__or2_1
X_05479_ _10224_/Q input64/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05479_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07218_ _07036_/A _07204_/B _07771_/B1 _10375_/Q vssd1 vssd1 vccd1 vccd1 _10375_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08198_ _08578_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _10934_/D sky130_fd_sc_hd__and2_1
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07149_ _10336_/Q _07145_/B _07188_/S _07040_/B vssd1 vssd1 vccd1 vccd1 _10336_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10160_ _11792_/Q _10176_/B vssd1 vssd1 vccd1 vccd1 _10160_/X sky130_fd_sc_hd__or2_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1006 input79/X vssd1 vssd1 vccd1 vccd1 _05751_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_105_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1017 _07021_/A vssd1 vssd1 vccd1 vccd1 _10105_/A1 sky130_fd_sc_hd__buf_6
X_10091_ _10182_/A0 _10087_/X _10090_/X _10155_/C1 vssd1 vssd1 vccd1 vccd1 _11747_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout1028 _10023_/A0 vssd1 vssd1 vccd1 vccd1 _10175_/A1 sky130_fd_sc_hd__buf_8
Xfanout1039 _08919_/A1 vssd1 vssd1 vccd1 vccd1 _09971_/A0 sky130_fd_sc_hd__clkbuf_8
XFILLER_134_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10993_ _11758_/CLK _10993_/D vssd1 vssd1 vccd1 vccd1 _10993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11614_ _11663_/CLK _11614_/D vssd1 vssd1 vccd1 vccd1 _11614_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_141_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11545_ _11801_/CLK _11545_/D vssd1 vssd1 vccd1 vccd1 _11545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11476_ _11477_/CLK _11476_/D vssd1 vssd1 vccd1 vccd1 _11476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10427_ _11284_/CLK _10427_/D vssd1 vssd1 vccd1 vccd1 _10427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ _11720_/CLK _10358_/D vssd1 vssd1 vccd1 vccd1 _10358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10289_ _10812_/CLK _10289_/D vssd1 vssd1 vccd1 vccd1 _10289_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06520_ _10665_/Q _09131_/A _06519_/X _06873_/D1 vssd1 vssd1 vccd1 vccd1 _06520_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06451_ _06535_/A _06450_/X _06449_/X _06664_/C1 vssd1 vssd1 vccd1 vccd1 _06451_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05402_ _10590_/Q _10589_/Q _05413_/S vssd1 vssd1 vccd1 vccd1 _05406_/A sky130_fd_sc_hd__mux2_1
X_09170_ _11429_/Q _09154_/X _09169_/X vssd1 vssd1 vccd1 vccd1 _11429_/D sky130_fd_sc_hd__a21o_1
X_06382_ _06900_/A _06353_/X _06364_/X _06381_/X vssd1 vssd1 vccd1 vccd1 _06382_/X
+ sky130_fd_sc_hd__a31o_1
X_08121_ _08578_/A _08121_/B vssd1 vssd1 vccd1 vccd1 _10887_/D sky130_fd_sc_hd__and2_1
X_05333_ _10847_/Q _10846_/Q _05394_/S vssd1 vssd1 vccd1 vccd1 _05334_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08052_ _08578_/A _08052_/B vssd1 vssd1 vccd1 vccd1 _10852_/D sky130_fd_sc_hd__and2_1
X_05264_ _05264_/A _05264_/B _05264_/C _05264_/D vssd1 vssd1 vccd1 vccd1 _05270_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07003_ _09540_/A _07003_/B vssd1 vssd1 vccd1 vccd1 _07003_/Y sky130_fd_sc_hd__nor2_2
XFILLER_31_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05195_ _06939_/A _11025_/Q vssd1 vssd1 vccd1 vccd1 _05195_/X sky130_fd_sc_hd__and2_1
XFILLER_116_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput109 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 _07042_/A sky130_fd_sc_hd__buf_6
X_08954_ _06945_/B _09540_/A _05472_/B _08953_/Y _05085_/Y vssd1 vssd1 vccd1 vccd1
+ _09830_/B sky130_fd_sc_hd__a2111o_4
XFILLER_9_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07905_ _10015_/A0 _10770_/Q _09218_/S vssd1 vssd1 vccd1 vccd1 _07906_/B sky130_fd_sc_hd__mux2_1
X_08885_ _08941_/A _08885_/B vssd1 vssd1 vccd1 vccd1 _11299_/D sky130_fd_sc_hd__or2_1
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07836_ _10047_/A1 _07839_/A2 _07961_/S _10731_/Q vssd1 vssd1 vccd1 vccd1 _10731_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07767_ _10687_/Q _07095_/X _07772_/S vssd1 vssd1 vccd1 vccd1 _10687_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09506_ _09492_/B _09528_/B _09504_/Y _09505_/X _09825_/A vssd1 vssd1 vccd1 vccd1
+ _11612_/D sky130_fd_sc_hd__o311a_1
X_06718_ _11331_/Q _09271_/A _06718_/B1 _11303_/Q _06718_/C1 vssd1 vssd1 vccd1 vccd1
+ _06718_/X sky130_fd_sc_hd__o221a_1
XFILLER_25_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07698_ _10646_/Q _07693_/Y _07697_/Y _08326_/B2 vssd1 vssd1 vccd1 vccd1 _10646_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06649_ _10348_/Q _06649_/A2 _06645_/X _06648_/X vssd1 vssd1 vccd1 vccd1 _06649_/X
+ sky130_fd_sc_hd__a211o_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _11590_/Q _11649_/Q _09440_/S vssd1 vssd1 vccd1 vccd1 _11590_/D sky130_fd_sc_hd__mux2_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09368_ _11542_/Q _09376_/B vssd1 vssd1 vccd1 vccd1 _09368_/X sky130_fd_sc_hd__or2_1
XFILLER_36_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08319_ _10080_/A0 _10998_/Q _08321_/S vssd1 vssd1 vccd1 vccd1 _10998_/D sky130_fd_sc_hd__mux2_1
XFILLER_138_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09299_ _09364_/A1 _09293_/X _09298_/X _09995_/C1 vssd1 vssd1 vccd1 vccd1 _11500_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_60 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 _05680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_82 _10213_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _11330_/CLK _11330_/D vssd1 vssd1 vccd1 vccd1 _11330_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_93 _09950_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11261_ _11262_/CLK _11261_/D vssd1 vssd1 vccd1 vccd1 _11261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10212_ _11808_/CLK _10212_/D vssd1 vssd1 vccd1 vccd1 _10212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11192_ _11251_/CLK _11192_/D vssd1 vssd1 vccd1 vccd1 _11192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10143_ _11784_/Q _10137_/X _10142_/X vssd1 vssd1 vccd1 vccd1 _11784_/D sky130_fd_sc_hd__a21o_1
XFILLER_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10074_ _10110_/A0 _11734_/Q _10082_/S vssd1 vssd1 vccd1 vccd1 _11734_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _11307_/CLK _10976_/D vssd1 vssd1 vccd1 vccd1 _10976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11528_ _11765_/CLK _11528_/D vssd1 vssd1 vccd1 vccd1 _11528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11459_ _11473_/CLK _11459_/D vssd1 vssd1 vccd1 vccd1 _11459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05951_ _06450_/A _10225_/Q vssd1 vssd1 vccd1 vccd1 _05951_/Y sky130_fd_sc_hd__nand2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08670_ _08670_/A _08670_/B vssd1 vssd1 vccd1 vccd1 _11189_/D sky130_fd_sc_hd__or2_1
XFILLER_61_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05882_ _06633_/A _05875_/X _05880_/X _06619_/A1 _05870_/X vssd1 vssd1 vccd1 vccd1
+ _05882_/X sky130_fd_sc_hd__o311a_1
XFILLER_94_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07621_ _09229_/A _08035_/S _07335_/X vssd1 vssd1 vccd1 vccd1 _07621_/X sky130_fd_sc_hd__a21o_1
XFILLER_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07552_ _07916_/A _07552_/B vssd1 vssd1 vccd1 vccd1 _10559_/D sky130_fd_sc_hd__or2_1
XFILLER_59_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06503_ _10793_/Q _06540_/A2 _06540_/B1 _10433_/Q vssd1 vssd1 vccd1 vccd1 _06503_/X
+ sky130_fd_sc_hd__o22a_1
X_07483_ _07076_/A _10520_/Q _07483_/S vssd1 vssd1 vccd1 vccd1 _07484_/B sky130_fd_sc_hd__mux2_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09222_ _09243_/B _07037_/B _09209_/Y _09221_/X vssd1 vssd1 vccd1 vccd1 _11460_/D
+ sky130_fd_sc_hd__a31o_1
X_06434_ _10705_/Q _09059_/A _09131_/A _10663_/Q _06433_/X vssd1 vssd1 vccd1 vccd1
+ _06434_/X sky130_fd_sc_hd__a221o_1
XFILLER_72_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09153_ _10158_/A _10136_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09171_/B sky130_fd_sc_hd__and3_4
X_06365_ _10753_/Q _06861_/B vssd1 vssd1 vccd1 vccd1 _06365_/X sky130_fd_sc_hd__or2_1
XFILLER_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08104_ _10876_/Q _08102_/S _07642_/S _07227_/B vssd1 vssd1 vccd1 vccd1 _10876_/D
+ sky130_fd_sc_hd__o22a_1
X_05316_ _10876_/Q _10875_/Q _05396_/S vssd1 vssd1 vccd1 vccd1 _05318_/C sky130_fd_sc_hd__mux2_1
X_09084_ _09111_/A1 _09082_/X _09083_/X _09092_/C1 vssd1 vssd1 vccd1 vccd1 _11389_/D
+ sky130_fd_sc_hd__o211a_1
X_06296_ _11526_/Q _09326_/A _09132_/A _11790_/Q _06295_/X vssd1 vssd1 vccd1 vccd1
+ _06296_/X sky130_fd_sc_hd__o221a_1
X_08035_ _09234_/A0 _10842_/Q _08035_/S vssd1 vssd1 vccd1 vccd1 _08036_/B sky130_fd_sc_hd__mux2_1
X_05247_ _05247_/A _05247_/B _05247_/C _05247_/D vssd1 vssd1 vccd1 vccd1 _05248_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput80 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__clkbuf_2
Xinput91 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__buf_2
XFILLER_116_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05178_ _05178_/A _05178_/B _05178_/C _05178_/D vssd1 vssd1 vccd1 vccd1 _05179_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_107_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09986_ _11680_/Q _09994_/B vssd1 vssd1 vccd1 vccd1 _09986_/X sky130_fd_sc_hd__or2_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08937_ _08937_/A1 _08940_/S _08936_/X _08937_/C1 vssd1 vssd1 vccd1 vccd1 _11327_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08868_ _09285_/A1 _11291_/Q _08874_/S vssd1 vssd1 vccd1 vccd1 _08869_/B sky130_fd_sc_hd__mux2_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07819_ _07819_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _07819_/Y sky130_fd_sc_hd__nor2_8
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08799_ _09216_/A0 _08802_/S _08798_/X _08921_/C1 vssd1 vssd1 vccd1 vccd1 _11255_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10830_ _11604_/CLK _10830_/D vssd1 vssd1 vccd1 vccd1 _10830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10761_ _11457_/CLK _10761_/D vssd1 vssd1 vccd1 vccd1 _10761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10692_ _11477_/CLK _10692_/D vssd1 vssd1 vccd1 vccd1 _10692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11313_ _11411_/CLK _11313_/D vssd1 vssd1 vccd1 vccd1 _11313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11244_ _11291_/CLK _11244_/D vssd1 vssd1 vccd1 vccd1 _11244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11175_ _11766_/CLK _11175_/D vssd1 vssd1 vccd1 vccd1 _11175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10126_ _07015_/A _11772_/Q _10134_/S vssd1 vssd1 vccd1 vccd1 _11772_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10057_ _11720_/Q _07143_/A _10057_/S vssd1 vssd1 vccd1 vccd1 _10058_/B sky130_fd_sc_hd__mux2_1
XFILLER_36_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10959_ _11683_/CLK _10959_/D vssd1 vssd1 vccd1 vccd1 _10959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11758_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_06150_ _10844_/Q _06643_/A2 _10010_/A _11137_/Q _06149_/X vssd1 vssd1 vccd1 vccd1
+ _06151_/C sky130_fd_sc_hd__o221a_1
XFILLER_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05101_ _09407_/A vssd1 vssd1 vccd1 vccd1 _05101_/Y sky130_fd_sc_hd__inv_2
X_06081_ _06450_/A _10226_/Q _06886_/A2 _06080_/X vssd1 vssd1 vccd1 vccd1 _10226_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_144_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout607 _05737_/X vssd1 vssd1 vccd1 vccd1 _06430_/A2 sky130_fd_sc_hd__clkbuf_8
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _11455_/Q _09877_/A2 _09874_/A2 _11451_/Q vssd1 vssd1 vccd1 vccd1 _09840_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout618 _06748_/A2 vssd1 vssd1 vccd1 vccd1 _07777_/A sky130_fd_sc_hd__buf_6
XFILLER_115_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout629 _05819_/B vssd1 vssd1 vccd1 vccd1 _06664_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_13__f_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_69_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09672_/B _09674_/A _09477_/A _09403_/Y vssd1 vssd1 vccd1 vccd1 _09771_/Y
+ sky130_fd_sc_hd__a211oi_4
X_06983_ _10259_/Q _06995_/B vssd1 vssd1 vccd1 vccd1 _06983_/X sky130_fd_sc_hd__or2_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08722_ _08810_/A _08722_/B vssd1 vssd1 vccd1 vccd1 _11217_/D sky130_fd_sc_hd__or2_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05934_ _06431_/A _05934_/B _05934_/C vssd1 vssd1 vccd1 vccd1 _05934_/X sky130_fd_sc_hd__or3_2
XFILLER_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05865_ _11767_/Q _05865_/B vssd1 vssd1 vccd1 vccd1 _05865_/X sky130_fd_sc_hd__or2_1
X_08653_ _11182_/Q _08437_/A _08748_/S _08303_/A vssd1 vssd1 vccd1 vccd1 _08653_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_96_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07604_ _10584_/Q _07598_/Y _07599_/Y _07013_/X vssd1 vssd1 vccd1 vccd1 _10584_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_96_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05796_ _10742_/Q _10009_/A _07819_/A _10300_/Q _05795_/X vssd1 vssd1 vccd1 vccd1
+ _05796_/X sky130_fd_sc_hd__o221a_1
X_08584_ _09396_/A0 _08589_/S _08583_/X _08831_/C1 vssd1 vssd1 vccd1 vccd1 _11147_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07535_ _07143_/A _10552_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _07536_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07466_ _07476_/A _07466_/B vssd1 vssd1 vccd1 vccd1 _10510_/D sky130_fd_sc_hd__or2_1
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09205_ _09214_/B _09208_/B vssd1 vssd1 vccd1 vccd1 _09205_/Y sky130_fd_sc_hd__nor2_4
X_06417_ _10943_/Q _06459_/A2 _06459_/B1 _11019_/Q vssd1 vssd1 vccd1 vccd1 _06417_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07397_ _07002_/A _10475_/Q _07429_/S vssd1 vssd1 vccd1 vccd1 _07398_/B sky130_fd_sc_hd__mux2_1
XFILLER_33_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09136_ _11413_/Q _09132_/X _09135_/X vssd1 vssd1 vccd1 vccd1 _11413_/D sky130_fd_sc_hd__a21o_1
X_06348_ _11567_/Q _09391_/A _09380_/A _11557_/Q vssd1 vssd1 vccd1 vccd1 _06348_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09067_ _09090_/A1 _09077_/B _08783_/A vssd1 vssd1 vccd1 vccd1 _09067_/X sky130_fd_sc_hd__a21o_1
X_06279_ _11694_/Q _09998_/A _06924_/A _11741_/Q _06344_/C1 vssd1 vssd1 vccd1 vccd1
+ _06279_/X sky130_fd_sc_hd__o221a_1
XFILLER_2_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08018_ _08469_/A _08011_/S _08017_/X _08841_/C1 vssd1 vssd1 vccd1 vccd1 _10833_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09969_ _10112_/A0 _11669_/Q _09975_/S vssd1 vssd1 vccd1 vccd1 _11669_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10813_ _11776_/CLK _10813_/D vssd1 vssd1 vccd1 vccd1 _10813_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _11801_/CLK _11793_/D vssd1 vssd1 vccd1 vccd1 _11793_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10744_ _11220_/CLK _10744_/D vssd1 vssd1 vccd1 vccd1 _10744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10675_ _11439_/CLK _10675_/D vssd1 vssd1 vccd1 vccd1 _10675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11227_ _11629_/CLK _11227_/D vssd1 vssd1 vccd1 vccd1 _11227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11158_ _11332_/CLK _11158_/D vssd1 vssd1 vccd1 vccd1 _11158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10109_ _10181_/A0 _11756_/Q _10118_/S vssd1 vssd1 vccd1 vccd1 _11756_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11089_ _11607_/CLK _11089_/D vssd1 vssd1 vccd1 vccd1 _11089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05650_ _11302_/Q _05543_/Y _05615_/Y _11298_/Q vssd1 vssd1 vccd1 vccd1 _05650_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05581_ _09552_/A1 _11387_/Q _11381_/Q _05078_/A vssd1 vssd1 vccd1 vccd1 _05581_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07320_ _08286_/A _08471_/B _10136_/C vssd1 vssd1 vccd1 vccd1 _08164_/B sky130_fd_sc_hd__and3_4
XFILLER_20_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07251_ _07036_/A _07665_/S _10058_/A vssd1 vssd1 vccd1 vccd1 _07251_/X sky130_fd_sc_hd__a21o_1
XFILLER_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06202_ _11109_/Q _06716_/A2 _06221_/A2 _11158_/Q vssd1 vssd1 vccd1 vccd1 _06202_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07182_ _10051_/A1 _10352_/Q _09243_/C vssd1 vssd1 vccd1 vccd1 _07183_/B sky130_fd_sc_hd__mux2_1
XFILLER_34_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06133_ _10940_/Q _06630_/A2 _06459_/B1 _11016_/Q vssd1 vssd1 vccd1 vccd1 _06133_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06064_ _11307_/Q _10009_/A _06060_/X _06063_/X vssd1 vssd1 vccd1 vccd1 _06064_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout404 _05401_/Y vssd1 vssd1 vccd1 vccd1 _09572_/C sky130_fd_sc_hd__buf_6
XFILLER_28_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout415 _05346_/Y vssd1 vssd1 vccd1 vccd1 _09567_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout426 _05281_/Y vssd1 vssd1 vccd1 vccd1 _09572_/B sky130_fd_sc_hd__buf_8
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout437 _05224_/Y vssd1 vssd1 vccd1 vccd1 _09873_/B1 sky130_fd_sc_hd__buf_4
X_09823_ _09823_/A _09823_/B vssd1 vssd1 vccd1 vccd1 _09823_/Y sky130_fd_sc_hd__xnor2_2
Xfanout448 _05157_/Y vssd1 vssd1 vccd1 vccd1 _09947_/A2 sky130_fd_sc_hd__buf_8
XFILLER_150_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout459 _08821_/A vssd1 vssd1 vccd1 vccd1 _08578_/A sky130_fd_sc_hd__buf_4
XFILLER_154_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09754_ _10539_/Q _09876_/B1 _09877_/B1 _10499_/Q _09753_/X vssd1 vssd1 vccd1 vccd1
+ _09757_/C sky130_fd_sc_hd__a221o_1
X_06966_ _10220_/Q _06965_/X _09416_/A vssd1 vssd1 vccd1 vccd1 _10220_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08705_ _11207_/Q _08705_/B vssd1 vssd1 vccd1 vccd1 _08705_/X sky130_fd_sc_hd__or2_1
X_05917_ _10770_/Q _06862_/A2 _05913_/X _05916_/X vssd1 vssd1 vccd1 vccd1 _05917_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_27_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09685_ _09703_/A _09685_/B vssd1 vssd1 vccd1 vccd1 _11635_/D sky130_fd_sc_hd__or2_1
X_06897_ _07689_/A _07689_/B vssd1 vssd1 vccd1 vccd1 _10180_/C sky130_fd_sc_hd__nand2_8
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _07005_/A _08637_/C _08635_/X vssd1 vssd1 vccd1 vccd1 _11172_/D sky130_fd_sc_hd__a21o_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05848_ _10682_/Q _06799_/A2 _05844_/X _05847_/X vssd1 vssd1 vccd1 vccd1 _05848_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08567_ _11138_/Q _07018_/A _08567_/S vssd1 vssd1 vccd1 vccd1 _08568_/B sky130_fd_sc_hd__mux2_1
X_05779_ _10364_/Q _07202_/A _05775_/X _05778_/X vssd1 vssd1 vccd1 vccd1 _05779_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07518_ _07930_/A _07518_/B vssd1 vssd1 vccd1 vccd1 _10543_/D sky130_fd_sc_hd__or2_1
XFILLER_80_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08498_ _08833_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _11099_/D sky130_fd_sc_hd__or2_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07449_ _07031_/A _07537_/B _07441_/Y _10501_/Q _09192_/A vssd1 vssd1 vccd1 vccd1
+ _10501_/D sky130_fd_sc_hd__a221o_1
XFILLER_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10460_ _11308_/CLK _10460_/D vssd1 vssd1 vccd1 vccd1 _10460_/Q sky130_fd_sc_hd__dfxtp_1
X_09119_ _09280_/A1 _09127_/B _09129_/B1 vssd1 vssd1 vccd1 vccd1 _09119_/X sky130_fd_sc_hd__a21o_1
X_10391_ _11743_/CLK _10391_/D vssd1 vssd1 vccd1 vccd1 _10391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11012_ _11733_/CLK _11012_/D vssd1 vssd1 vccd1 vccd1 _11012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout960 input92/X vssd1 vssd1 vccd1 vccd1 _08661_/A sky130_fd_sc_hd__clkbuf_16
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout971 input90/X vssd1 vssd1 vccd1 vccd1 _08931_/A1 sky130_fd_sc_hd__clkbuf_16
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout982 _08669_/A0 vssd1 vssd1 vccd1 vccd1 _07303_/A sky130_fd_sc_hd__clkbuf_16
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 _07690_/B vssd1 vssd1 vccd1 vccd1 _06392_/C1 sky130_fd_sc_hd__buf_4
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1084 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1084/HI io_oeb[14] sky130_fd_sc_hd__conb_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1095 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1095/HI io_oeb[25] sky130_fd_sc_hd__conb_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _11776_/CLK _11776_/D vssd1 vssd1 vccd1 vccd1 _11776_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10727_ _10727_/CLK _10727_/D vssd1 vssd1 vccd1 vccd1 _10727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10658_ _10666_/CLK _10658_/D vssd1 vssd1 vccd1 vccd1 _10658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10589_ _11280_/CLK _10589_/D vssd1 vssd1 vccd1 vccd1 _10589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06820_ _10530_/Q _06873_/A2 _06710_/B _10735_/Q _06819_/X vssd1 vssd1 vccd1 vccd1
+ _06820_/X sky130_fd_sc_hd__o221a_1
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06751_ _10350_/Q _06766_/A2 _06750_/X _06878_/C1 vssd1 vssd1 vccd1 vccd1 _06751_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05702_ _11118_/Q _05561_/Y _05585_/Y _11117_/Q _05701_/X vssd1 vssd1 vccd1 vccd1
+ _05703_/C sky130_fd_sc_hd__a221o_1
X_06682_ _06577_/A _10238_/Q _06855_/B vssd1 vssd1 vccd1 vccd1 _06682_/X sky130_fd_sc_hd__a21o_1
X_09470_ _09475_/A _09470_/B vssd1 vssd1 vccd1 vccd1 _09470_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08421_ _08893_/A1 _08404_/S _08420_/X _08919_/C1 vssd1 vssd1 vccd1 vccd1 _11051_/D
+ sky130_fd_sc_hd__o211a_1
X_05633_ _05633_/A _05633_/B vssd1 vssd1 vccd1 vccd1 _05633_/Y sky130_fd_sc_hd__nor2_8
XFILLER_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05564_ _11795_/Q _05618_/A1 _05620_/B2 _11793_/Q _05562_/X vssd1 vssd1 vccd1 vccd1
+ _05567_/A sky130_fd_sc_hd__a221o_4
Xclkbuf_leaf_53_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11235_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08352_ _11019_/Q _08362_/B vssd1 vssd1 vccd1 vccd1 _08352_/X sky130_fd_sc_hd__or2_1
XFILLER_71_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07303_ _07303_/A _07613_/A vssd1 vssd1 vccd1 vccd1 _07303_/X sky130_fd_sc_hd__or2_4
X_05495_ _10240_/Q input51/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05495_/X sky130_fd_sc_hd__mux2_1
X_08283_ _08893_/A1 _08245_/X _08282_/X _09092_/C1 vssd1 vssd1 vccd1 vccd1 _10973_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07234_ _07108_/X _10385_/Q _07246_/S vssd1 vssd1 vccd1 vccd1 _10385_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07165_ _07790_/A _07165_/B vssd1 vssd1 vccd1 vccd1 _10343_/D sky130_fd_sc_hd__or2_1
XFILLER_117_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06116_ _11318_/Q _09271_/A _06718_/B1 _11290_/Q _06718_/C1 vssd1 vssd1 vccd1 vccd1
+ _06119_/A sky130_fd_sc_hd__o221a_1
XFILLER_145_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07096_ _10303_/Q _07095_/X _07109_/S vssd1 vssd1 vccd1 vccd1 _10303_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06047_ _10342_/Q _07152_/A _06046_/X _06651_/C1 vssd1 vssd1 vccd1 vccd1 _06047_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout212 _07959_/S vssd1 vssd1 vccd1 vccd1 _07821_/A sky130_fd_sc_hd__buf_6
XFILLER_114_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout223 _07233_/S vssd1 vssd1 vccd1 vccd1 _07249_/S sky130_fd_sc_hd__buf_8
XFILLER_8_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout234 _07044_/S vssd1 vssd1 vccd1 vccd1 _07038_/S sky130_fd_sc_hd__buf_8
Xfanout245 _08907_/X vssd1 vssd1 vccd1 vccd1 _08945_/A2 sky130_fd_sc_hd__buf_6
Xfanout256 _08650_/X vssd1 vssd1 vccd1 vccd1 _08742_/S sky130_fd_sc_hd__clkbuf_4
X_09806_ _10282_/Q _09566_/C _09572_/C _10530_/Q vssd1 vssd1 vccd1 vccd1 _09806_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout267 _08832_/S vssd1 vssd1 vccd1 vccd1 _08838_/S sky130_fd_sc_hd__buf_6
Xfanout278 _07994_/X vssd1 vssd1 vccd1 vccd1 _08011_/S sky130_fd_sc_hd__buf_6
XFILLER_75_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout289 _07853_/Y vssd1 vssd1 vccd1 vccd1 _07893_/B sky130_fd_sc_hd__buf_4
X_07998_ _08833_/A _07998_/B vssd1 vssd1 vccd1 vccd1 _10823_/D sky130_fd_sc_hd__or2_1
XFILLER_41_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09737_ _10338_/Q _09874_/A2 _09565_/D _10349_/Q vssd1 vssd1 vccd1 vccd1 _09737_/X
+ sky130_fd_sc_hd__a22o_1
X_06949_ _09538_/B input6/X _08955_/A vssd1 vssd1 vccd1 vccd1 _06950_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09668_ _09668_/A _09668_/B _09668_/C _09668_/D vssd1 vssd1 vccd1 vccd1 _09669_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _08846_/A0 _11164_/Q _08621_/S vssd1 vssd1 vccd1 vccd1 _08620_/B sky130_fd_sc_hd__mux2_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09827_/A _09823_/B _09823_/A vssd1 vssd1 vccd1 vccd1 _09599_/X sky130_fd_sc_hd__or3b_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11702_/CLK _11630_/D vssd1 vssd1 vccd1 vccd1 _11630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11561_ _11675_/CLK _11561_/D vssd1 vssd1 vccd1 vccd1 _11561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10512_ _11698_/CLK _10512_/D vssd1 vssd1 vccd1 vccd1 _10512_/Q sky130_fd_sc_hd__dfxtp_1
X_11492_ _11497_/CLK _11492_/D vssd1 vssd1 vccd1 vccd1 _11492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10443_ _11768_/CLK _10443_/D vssd1 vssd1 vccd1 vccd1 _10443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10374_ _11713_/CLK _10374_/D vssd1 vssd1 vccd1 vccd1 _10374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout790 _06737_/B1 vssd1 vssd1 vccd1 vccd1 _08972_/A sky130_fd_sc_hd__buf_8
XFILLER_24_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_150 _06789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _07617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 _10013_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_194 _07021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11759_ _11765_/CLK _11759_/D vssd1 vssd1 vccd1 vccd1 _11759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05280_ _05280_/A _05280_/B _05280_/C _05280_/D vssd1 vssd1 vccd1 vccd1 _05281_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_140_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08970_ _11338_/Q _08970_/A1 _08970_/S vssd1 vssd1 vccd1 vccd1 _11338_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_100_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _10808_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07921_ _09182_/A0 _10778_/Q _09218_/S vssd1 vssd1 vccd1 vccd1 _07922_/B sky130_fd_sc_hd__mux2_1
XFILLER_151_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07852_ _08901_/A1 _10745_/Q _07852_/S vssd1 vssd1 vccd1 vccd1 _10745_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06803_ _10493_/Q _06803_/A2 _06799_/X _06802_/X vssd1 vssd1 vccd1 vccd1 _06803_/X
+ sky130_fd_sc_hd__o211a_2
Xinput1 io_in[5] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_151_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07783_ _10015_/A0 _10699_/Q _07817_/S vssd1 vssd1 vccd1 vccd1 _07784_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09522_ _09525_/A _09522_/B _09522_/C _09528_/B vssd1 vssd1 vccd1 vccd1 _09523_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06734_ _06878_/C1 _06732_/X _06733_/X _06743_/B vssd1 vssd1 vccd1 vccd1 _06734_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09453_ _05372_/S _09475_/A _09452_/Y _09407_/A vssd1 vssd1 vccd1 vccd1 _11596_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06665_ _11615_/Q _06665_/A2 _06663_/X _06853_/A3 _06664_/X vssd1 vssd1 vccd1 vccd1
+ _10237_/D sky130_fd_sc_hd__a221o_1
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08404_ _08876_/A0 _11043_/Q _08404_/S vssd1 vssd1 vccd1 vccd1 _08405_/B sky130_fd_sc_hd__mux2_1
X_05616_ _05616_/A1 _11376_/Q _11373_/Q _11626_/Q vssd1 vssd1 vccd1 vccd1 _05616_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09384_ _09395_/A0 _11551_/Q _09390_/S vssd1 vssd1 vccd1 vccd1 _11551_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06596_ _10820_/Q _06639_/B1 _08469_/B _11085_/Q vssd1 vssd1 vccd1 vccd1 _06596_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_71_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08335_ _11010_/Q _08323_/Y _08324_/Y _07335_/X vssd1 vssd1 vccd1 vccd1 _11010_/D
+ sky130_fd_sc_hd__o22a_1
X_05547_ _05619_/A1 _11497_/Q _11493_/Q _05619_/B2 _05545_/X vssd1 vssd1 vccd1 vccd1
+ _05547_/X sky130_fd_sc_hd__a221o_1
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05478_ _10223_/Q input53/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05478_/X sky130_fd_sc_hd__mux2_1
X_08266_ _08876_/A0 _10965_/Q _08276_/S vssd1 vssd1 vccd1 vccd1 _08267_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07217_ _07143_/A _07204_/B _07771_/B1 _10374_/Q vssd1 vssd1 vccd1 vccd1 _10374_/D
+ sky130_fd_sc_hd__a22o_1
X_08197_ _10934_/Q _10135_/A0 _08197_/S vssd1 vssd1 vccd1 vccd1 _08198_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07148_ _10335_/Q _07150_/A2 _07188_/S _07451_/B vssd1 vssd1 vccd1 vccd1 _10335_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07079_ _07036_/A _07074_/S _07078_/X _07141_/B vssd1 vssd1 vccd1 vccd1 _10298_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10090_ _11747_/Q _10104_/B vssd1 vssd1 vccd1 vccd1 _10090_/X sky130_fd_sc_hd__or2_1
Xfanout1007 _10190_/A0 vssd1 vssd1 vccd1 vccd1 _10118_/A0 sky130_fd_sc_hd__buf_4
Xfanout1018 _10177_/A1 vssd1 vssd1 vccd1 vccd1 _07021_/A sky130_fd_sc_hd__buf_12
XFILLER_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1029 input115/X vssd1 vssd1 vccd1 vccd1 _10023_/A0 sky130_fd_sc_hd__buf_12
XFILLER_0_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10992_ _11763_/CLK _10992_/D vssd1 vssd1 vccd1 vccd1 _10992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11812_/CLK _11613_/D vssd1 vssd1 vccd1 vccd1 _11613_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11544_ _11684_/CLK _11544_/D vssd1 vssd1 vccd1 vccd1 _11544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11475_ _11745_/CLK _11475_/D vssd1 vssd1 vccd1 vccd1 _11475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10426_ _11233_/CLK _10426_/D vssd1 vssd1 vccd1 vccd1 _10426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10357_ _10727_/CLK _10357_/D vssd1 vssd1 vccd1 vccd1 _10357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _11710_/CLK _10288_/D vssd1 vssd1 vccd1 vccd1 _10288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06450_ _06450_/A _10232_/Q vssd1 vssd1 vccd1 vccd1 _06450_/X sky130_fd_sc_hd__and2_1
XFILLER_34_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05401_ _05401_/A _05401_/B vssd1 vssd1 vccd1 vccd1 _05401_/Y sky130_fd_sc_hd__nor2_8
X_06381_ _06743_/B _06375_/X _06380_/X _07081_/A vssd1 vssd1 vccd1 vccd1 _06381_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08120_ _10887_/Q _10135_/A0 _08120_/S vssd1 vssd1 vccd1 vccd1 _08121_/B sky130_fd_sc_hd__mux2_1
X_05332_ _10852_/Q _10851_/Q _05399_/S vssd1 vssd1 vccd1 vccd1 _05334_/C sky130_fd_sc_hd__mux2_1
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05263_ _10438_/Q _10437_/Q _05396_/S vssd1 vssd1 vccd1 vccd1 _05264_/D sky130_fd_sc_hd__mux2_1
X_08051_ _10852_/Q _10135_/A0 _08051_/S vssd1 vssd1 vccd1 vccd1 _08052_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07002_ _07002_/A _07107_/B vssd1 vssd1 vccd1 vccd1 _07225_/A sky130_fd_sc_hd__and2_2
XFILLER_127_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05194_ _05419_/S _11068_/Q vssd1 vssd1 vccd1 vccd1 _05194_/X sky130_fd_sc_hd__and2b_1
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08953_ _05300_/S _08956_/B _09540_/A vssd1 vssd1 vccd1 vccd1 _08953_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07904_ _07904_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07904_/X sky130_fd_sc_hd__or2_1
XFILLER_9_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08884_ _08937_/A1 _11299_/Q _08884_/S vssd1 vssd1 vccd1 vccd1 _08885_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07835_ _07031_/A _07839_/A2 _07959_/S _10730_/Q vssd1 vssd1 vccd1 vccd1 _10730_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07766_ _10686_/Q _07617_/X _07772_/S vssd1 vssd1 vccd1 vccd1 _10686_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09505_ _09525_/A _09522_/B _09504_/B _09489_/C _11612_/Q vssd1 vssd1 vccd1 vccd1
+ _09505_/X sky130_fd_sc_hd__a41o_1
X_06717_ _11051_/Q _06735_/A2 _06717_/B1 _10973_/Q _06716_/X vssd1 vssd1 vccd1 vccd1
+ _06720_/A sky130_fd_sc_hd__o221a_1
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07697_ _08439_/A _08589_/S vssd1 vssd1 vccd1 vccd1 _07697_/Y sky130_fd_sc_hd__nand2_2
XFILLER_13_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _11589_/Q _11648_/Q _09440_/S vssd1 vssd1 vccd1 vccd1 _11589_/D sky130_fd_sc_hd__mux2_1
X_06648_ _10757_/Q _06648_/A2 _06647_/X _06873_/D1 vssd1 vssd1 vccd1 vccd1 _06648_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09985_/A1 _09359_/X _09366_/X _10177_/C1 vssd1 vssd1 vccd1 vccd1 _11541_/D
+ sky130_fd_sc_hd__o211a_1
X_06579_ _11613_/Q _05819_/Y _06577_/X _06622_/B2 _06578_/X vssd1 vssd1 vccd1 vccd1
+ _10235_/D sky130_fd_sc_hd__a221o_1
XFILLER_21_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08318_ _10115_/A0 _10997_/Q _08321_/S vssd1 vssd1 vccd1 vccd1 _10997_/D sky130_fd_sc_hd__mux2_1
X_09298_ _11500_/Q _09310_/B vssd1 vssd1 vccd1 vccd1 _09298_/X sky130_fd_sc_hd__or2_1
XANTENNA_50 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 _05704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_83 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ _09114_/A1 _08276_/S _08248_/X _09092_/C1 vssd1 vssd1 vccd1 vccd1 _10956_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_94 _09950_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11260_ _11262_/CLK _11260_/D vssd1 vssd1 vccd1 vccd1 _11260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10211_ _11811_/CLK _10211_/D vssd1 vssd1 vccd1 vccd1 _10211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11191_ _11251_/CLK _11191_/D vssd1 vssd1 vccd1 vccd1 _11191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10142_ _10142_/A1 _10154_/B _10156_/B1 vssd1 vssd1 vccd1 vccd1 _10142_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput190 _05496_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_4
X_10073_ _10181_/A0 _11733_/Q _10082_/S vssd1 vssd1 vccd1 vccd1 _11733_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10975_ _11307_/CLK _10975_/D vssd1 vssd1 vccd1 vccd1 _10975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11527_ _11527_/CLK _11527_/D vssd1 vssd1 vccd1 vccd1 _11527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11458_ _11458_/CLK _11458_/D vssd1 vssd1 vccd1 vccd1 _11458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10409_ _10782_/CLK _10409_/D vssd1 vssd1 vccd1 vccd1 _10409_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_3_4_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11389_ _11393_/CLK _11389_/D vssd1 vssd1 vccd1 vccd1 _11389_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_12__f_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_88_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_97_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05950_ _05950_/A _05950_/B vssd1 vssd1 vccd1 vccd1 _10224_/D sky130_fd_sc_hd__or2_1
XFILLER_87_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05881_ _07151_/B _05854_/X _05859_/X _05843_/X vssd1 vssd1 vccd1 vccd1 _05881_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_27_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07620_ _10595_/Q _07613_/Y _07614_/Y _07333_/X vssd1 vssd1 vccd1 vccd1 _10595_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07551_ _10019_/A0 _10559_/Q _07589_/S vssd1 vssd1 vccd1 vccd1 _07552_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06502_ _11281_/Q _06539_/A2 _06539_/B1 _10595_/Q _06624_/C1 vssd1 vssd1 vccd1 vccd1
+ _06502_/X sky130_fd_sc_hd__o221a_2
X_07482_ _10043_/A _07482_/B vssd1 vssd1 vccd1 vccd1 _10519_/D sky130_fd_sc_hd__or2_1
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ _11460_/Q _09243_/B _09221_/C vssd1 vssd1 vccd1 vccd1 _09221_/X sky130_fd_sc_hd__and3_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06433_ _10345_/Q _06649_/A2 _08971_/A _10564_/Q vssd1 vssd1 vccd1 vccd1 _06433_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ _11421_/Q _09132_/X _09151_/X vssd1 vssd1 vccd1 vccd1 _11421_/D sky130_fd_sc_hd__a21o_1
XFILLER_124_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06364_ _07297_/A _06364_/B _06364_/C vssd1 vssd1 vccd1 vccd1 _06364_/X sky130_fd_sc_hd__or3_2
X_08103_ _08819_/A _08103_/B vssd1 vssd1 vccd1 vccd1 _10875_/D sky130_fd_sc_hd__or2_1
X_05315_ _10880_/Q _10879_/Q _05392_/S vssd1 vssd1 vccd1 vccd1 _05318_/B sky130_fd_sc_hd__mux2_1
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06295_ _11800_/Q _10159_/A _09293_/A _11506_/Q vssd1 vssd1 vccd1 vccd1 _06295_/X
+ sky130_fd_sc_hd__o22a_1
X_09083_ _11389_/Q _09099_/B vssd1 vssd1 vccd1 vccd1 _09083_/X sky130_fd_sc_hd__or2_1
X_08034_ _08789_/A1 _08035_/S _08033_/X _07011_/B vssd1 vssd1 vccd1 vccd1 _10841_/D
+ sky130_fd_sc_hd__o211a_1
Xinput70 wb_rom_val[6] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_2
X_05246_ _10868_/Q _10867_/Q _06942_/A vssd1 vssd1 vccd1 vccd1 _05247_/D sky130_fd_sc_hd__mux2_1
Xinput81 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput92 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__buf_8
XFILLER_116_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05177_ _11182_/Q _11181_/Q _05427_/S vssd1 vssd1 vccd1 vccd1 _05178_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09985_ _09985_/A1 _09977_/X _09984_/X _09995_/C1 vssd1 vssd1 vccd1 vccd1 _11679_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08936_ _11327_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08936_/X sky130_fd_sc_hd__or2_1
XFILLER_131_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08867_ _08869_/A _08867_/B vssd1 vssd1 vccd1 vccd1 _11290_/D sky130_fd_sc_hd__or2_1
XFILLER_40_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07818_ _07818_/A _07818_/B vssd1 vssd1 vccd1 vccd1 _10716_/D sky130_fd_sc_hd__or2_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08798_ _11255_/Q _08804_/B vssd1 vssd1 vccd1 vccd1 _08798_/X sky130_fd_sc_hd__or2_1
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11652_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07749_ _07933_/A0 _07755_/A2 _07748_/X _07902_/C1 vssd1 vssd1 vccd1 vccd1 _10675_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10760_ _10808_/CLK _10760_/D vssd1 vssd1 vccd1 vccd1 _10760_/Q sky130_fd_sc_hd__dfxtp_1
X_09419_ _11649_/Q _11578_/Q _09704_/B vssd1 vssd1 vccd1 vccd1 _11578_/D sky130_fd_sc_hd__mux2_1
X_10691_ _10725_/CLK _10691_/D vssd1 vssd1 vccd1 vccd1 _10691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ _11312_/CLK _11312_/D vssd1 vssd1 vccd1 vccd1 _11312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11243_ _11243_/CLK _11243_/D vssd1 vssd1 vccd1 vccd1 _11243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11174_ _11269_/CLK _11174_/D vssd1 vssd1 vccd1 vccd1 _11174_/Q sky130_fd_sc_hd__dfxtp_1
X_10125_ _07052_/A _11771_/Q _10134_/S vssd1 vssd1 vccd1 vccd1 _11771_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10056_ _10056_/A _10056_/B vssd1 vssd1 vccd1 vccd1 _11719_/D sky130_fd_sc_hd__or2_1
XFILLER_87_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10958_ _11243_/CLK _10958_/D vssd1 vssd1 vccd1 vccd1 _10958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10889_ _10939_/CLK _10889_/D vssd1 vssd1 vccd1 vccd1 _10889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05100_ _10215_/Q input74/X vssd1 vssd1 vccd1 vccd1 _05100_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06080_ _05692_/X _06622_/A2 _06078_/X _06079_/Y vssd1 vssd1 vccd1 vccd1 _06080_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_78_wb_clk_i clkbuf_leaf_85_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11332_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout608 _06228_/A2 vssd1 vssd1 vccd1 vccd1 _07994_/A sky130_fd_sc_hd__buf_6
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout619 _06748_/A2 vssd1 vssd1 vccd1 vccd1 _07778_/A sky130_fd_sc_hd__buf_6
XFILLER_63_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _11646_/Q _09769_/X _09770_/S vssd1 vssd1 vccd1 vccd1 _11646_/D sky130_fd_sc_hd__mux2_1
X_06982_ _10183_/A0 _06976_/X _06981_/X _06996_/C1 vssd1 vssd1 vccd1 vccd1 _10258_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _11217_/Q _10132_/A0 _08726_/S vssd1 vssd1 vccd1 vccd1 _08722_/B sky130_fd_sc_hd__mux2_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05933_ _10911_/Q _07046_/A _05929_/X _05932_/X vssd1 vssd1 vccd1 vccd1 _05934_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08652_ _07303_/X _08748_/S _08651_/X _08427_/A vssd1 vssd1 vccd1 vccd1 _11181_/D
+ sky130_fd_sc_hd__o211a_1
X_05864_ _05864_/A _05864_/B _05864_/C vssd1 vssd1 vccd1 vccd1 _05864_/X sky130_fd_sc_hd__and3_1
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07603_ _10583_/Q _07597_/Y _07600_/Y _07008_/X vssd1 vssd1 vccd1 vccd1 _10583_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08583_ _11147_/Q _08591_/B vssd1 vssd1 vccd1 vccd1 _08583_/X sky130_fd_sc_hd__or2_1
XFILLER_19_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05795_ _10435_/Q _06634_/B1 _07190_/A _10601_/Q vssd1 vssd1 vccd1 vccd1 _05795_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07534_ _07936_/A _07534_/B vssd1 vssd1 vccd1 vccd1 _10551_/D sky130_fd_sc_hd__or2_1
XFILLER_81_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07465_ _07057_/A _10510_/Q _07477_/S vssd1 vssd1 vccd1 vccd1 _07466_/B sky130_fd_sc_hd__mux2_1
X_09204_ _11450_/Q _09190_/Y _09193_/Y _07043_/X vssd1 vssd1 vccd1 vccd1 _11450_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06416_ _10652_/Q _06629_/A2 _06589_/A2 _11097_/Q _07690_/B vssd1 vssd1 vccd1 vccd1
+ _06416_/X sky130_fd_sc_hd__o221a_1
X_07396_ _10039_/A _07396_/B vssd1 vssd1 vccd1 vccd1 _10474_/D sky130_fd_sc_hd__or2_1
XFILLER_33_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09135_ _09275_/A1 _09149_/B _10166_/B1 vssd1 vssd1 vccd1 vccd1 _09135_/X sky130_fd_sc_hd__a21o_1
X_06347_ _11517_/Q _09314_/A _06343_/X _06346_/X vssd1 vssd1 vccd1 vccd1 _06353_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ _09276_/A1 _09060_/X _09065_/X _09078_/C1 vssd1 vssd1 vccd1 vccd1 _11381_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06278_ _11674_/Q _09965_/A _06284_/B1 _10999_/Q vssd1 vssd1 vccd1 vccd1 _06278_/X
+ sky130_fd_sc_hd__o22a_1
X_08017_ _10833_/Q _08091_/C vssd1 vssd1 vccd1 vccd1 _08017_/X sky130_fd_sc_hd__or2_1
X_05229_ _06967_/A _11002_/Q vssd1 vssd1 vccd1 vccd1 _05229_/X sky130_fd_sc_hd__and2_1
XFILLER_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09968_ _10111_/A0 _11668_/Q _09975_/S vssd1 vssd1 vccd1 vccd1 _11668_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08919_ _08919_/A1 _08945_/A2 _08918_/X _08919_/C1 vssd1 vssd1 vccd1 vccd1 _11318_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09899_ _09899_/A _09899_/B _09899_/C _09899_/D vssd1 vssd1 vccd1 vccd1 _09907_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_92_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _10812_/CLK _10812_/D vssd1 vssd1 vccd1 vccd1 _10812_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _11792_/CLK _11792_/D vssd1 vssd1 vccd1 vccd1 _11792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10743_ _11770_/CLK _10743_/D vssd1 vssd1 vccd1 vccd1 _10743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10674_ _11458_/CLK _10674_/D vssd1 vssd1 vccd1 vccd1 _10674_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11226_ _11651_/CLK _11226_/D vssd1 vssd1 vccd1 vccd1 _11226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11157_ _11251_/CLK _11157_/D vssd1 vssd1 vccd1 vccd1 _11157_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_136_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10108_ _10108_/A _10108_/B _10108_/C vssd1 vssd1 vccd1 vccd1 _10118_/S sky130_fd_sc_hd__or3_4
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11088_ _11312_/CLK _11088_/D vssd1 vssd1 vccd1 vccd1 _11088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10039_ _10039_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _11709_/D sky130_fd_sc_hd__or2_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_125_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11703_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_97_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05580_ _05616_/A1 _11386_/Q _11383_/Q _05077_/A vssd1 vssd1 vccd1 vccd1 _05580_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07250_ _07143_/X _07665_/S _07249_/S _10394_/Q _09214_/B vssd1 vssd1 vccd1 vccd1
+ _10394_/D sky130_fd_sc_hd__a221o_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06201_ _11195_/Q _06736_/A2 _06737_/B1 _10961_/Q vssd1 vssd1 vccd1 vccd1 _06201_/X
+ sky130_fd_sc_hd__o22a_1
X_07181_ _07918_/A _07181_/B vssd1 vssd1 vccd1 vccd1 _10351_/D sky130_fd_sc_hd__or2_1
XFILLER_30_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06132_ _10825_/Q _06415_/A2 _08300_/A _11270_/Q vssd1 vssd1 vccd1 vccd1 _06132_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06063_ _11223_/Q _06238_/A2 _06061_/X _06062_/X vssd1 vssd1 vccd1 vccd1 _06063_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout405 _05401_/Y vssd1 vssd1 vccd1 vccd1 _09886_/B1 sky130_fd_sc_hd__buf_4
XFILLER_113_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout416 _05335_/Y vssd1 vssd1 vccd1 vccd1 _09571_/C sky130_fd_sc_hd__buf_8
Xfanout427 _05281_/Y vssd1 vssd1 vccd1 vccd1 _09872_/A2 sky130_fd_sc_hd__buf_6
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09822_ _09825_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _11654_/D sky130_fd_sc_hd__and2_1
XFILLER_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout438 _05214_/Y vssd1 vssd1 vccd1 vccd1 _09566_/B sky130_fd_sc_hd__buf_8
XFILLER_28_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout449 _05157_/Y vssd1 vssd1 vccd1 vccd1 _09573_/A sky130_fd_sc_hd__buf_4
XFILLER_58_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09753_ _10553_/Q _09953_/B1 _09884_/A2 _10541_/Q vssd1 vssd1 vccd1 vccd1 _09753_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_100_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06965_ _11664_/Q _05474_/B _06964_/X vssd1 vssd1 vccd1 vccd1 _06965_/X sky130_fd_sc_hd__a21o_2
XFILLER_80_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08704_ _09237_/A0 _08695_/S _08703_/X _07003_/B vssd1 vssd1 vccd1 vccd1 _11206_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05916_ _10340_/Q _06766_/A2 _05915_/X _06808_/C1 vssd1 vssd1 vccd1 vccd1 _05916_/X
+ sky130_fd_sc_hd__o211a_1
X_09684_ _05426_/S _09682_/B _09682_/Y _11635_/Q _09683_/X vssd1 vssd1 vccd1 vccd1
+ _09685_/B sky130_fd_sc_hd__o221a_1
X_06896_ _07690_/A _07298_/B vssd1 vssd1 vccd1 vccd1 _09015_/B sky130_fd_sc_hd__nor2_2
XFILLER_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ _11172_/Q _08437_/A _08140_/S _08438_/A vssd1 vssd1 vccd1 vccd1 _08635_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05847_ _11697_/Q _06857_/B1 _05846_/X _06997_/A vssd1 vssd1 vccd1 vccd1 _05847_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _11137_/Q _08567_/S _08563_/Y _07095_/B vssd1 vssd1 vccd1 vccd1 _11137_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_1280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05778_ _11696_/Q _10009_/A _05777_/X _06997_/A vssd1 vssd1 vccd1 vccd1 _05778_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07517_ _09182_/A0 _10543_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _07518_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08497_ _07104_/A _11099_/Q _08497_/S vssd1 vssd1 vccd1 vccd1 _08498_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07448_ _07028_/A _07537_/B _07441_/Y _10500_/Q _09228_/A vssd1 vssd1 vccd1 vccd1
+ _10500_/D sky130_fd_sc_hd__a221o_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07379_ _10464_/Q _07393_/S _07655_/S _07229_/B vssd1 vssd1 vccd1 vccd1 _10464_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09118_ _11405_/Q _09110_/X _09117_/X vssd1 vssd1 vccd1 vccd1 _11405_/D sky130_fd_sc_hd__a21o_1
X_10390_ _11477_/CLK _10390_/D vssd1 vssd1 vccd1 vccd1 _10390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09049_ _09283_/A1 _09055_/B _09290_/B1 vssd1 vssd1 vccd1 vccd1 _09049_/X sky130_fd_sc_hd__a21o_1
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11011_ _11023_/CLK _11011_/D vssd1 vssd1 vccd1 vccd1 _11011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout950 input94/X vssd1 vssd1 vccd1 vccd1 _08939_/A1 sky130_fd_sc_hd__buf_8
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout961 _08935_/A1 vssd1 vssd1 vccd1 vccd1 _08883_/A1 sky130_fd_sc_hd__buf_6
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout972 input89/X vssd1 vssd1 vccd1 vccd1 _07059_/A sky130_fd_sc_hd__buf_12
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout983 input88/X vssd1 vssd1 vccd1 vccd1 _08669_/A0 sky130_fd_sc_hd__clkbuf_16
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 _07298_/B vssd1 vssd1 vccd1 vccd1 _07690_/B sky130_fd_sc_hd__buf_12
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1085 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1085/HI io_oeb[15] sky130_fd_sc_hd__conb_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1096 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1096/HI io_oeb[26] sky130_fd_sc_hd__conb_1
XFILLER_61_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11779_/CLK _11775_/D vssd1 vssd1 vccd1 vccd1 _11775_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _10727_/CLK _10726_/D vssd1 vssd1 vccd1 vccd1 _10726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10657_ _11644_/CLK _10657_/D vssd1 vssd1 vccd1 vccd1 _10657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10588_ _11280_/CLK _10588_/D vssd1 vssd1 vccd1 vccd1 _10588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11209_ _11770_/CLK _11209_/D vssd1 vssd1 vccd1 vccd1 _11209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06750_ _10783_/Q _06875_/A2 _06875_/B1 _10673_/Q _06749_/X vssd1 vssd1 vccd1 vccd1
+ _06750_/X sky130_fd_sc_hd__o221a_1
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05701_ _11119_/Q _05579_/Y _05597_/Y _11110_/Q vssd1 vssd1 vccd1 vccd1 _05701_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06681_ _11168_/Q _06735_/B1 _06678_/X _06680_/X vssd1 vssd1 vccd1 vccd1 _06681_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_63_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08420_ _11051_/Q _08422_/B vssd1 vssd1 vccd1 vccd1 _08420_/X sky130_fd_sc_hd__or2_1
X_05632_ _11788_/Q _11627_/Q _05079_/A _11782_/Q _05631_/X vssd1 vssd1 vccd1 vccd1
+ _05633_/B sky130_fd_sc_hd__a221o_4
XFILLER_149_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08351_ _10190_/A0 _08360_/S _08350_/X _08351_/C1 vssd1 vssd1 vccd1 vccd1 _11018_/D
+ sky130_fd_sc_hd__o211a_1
X_05563_ _11800_/Q _09552_/A1 _05078_/A _11794_/Q vssd1 vssd1 vccd1 vccd1 _05563_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07302_ _08323_/A _08760_/S vssd1 vssd1 vccd1 vccd1 _07302_/Y sky130_fd_sc_hd__nand2_2
XFILLER_71_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08282_ _10973_/Q _08284_/B vssd1 vssd1 vccd1 vccd1 _08282_/X sky130_fd_sc_hd__or2_1
X_05494_ _10239_/Q input50/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05494_/X sky130_fd_sc_hd__mux2_1
X_07233_ _07232_/X _10384_/Q _07233_/S vssd1 vssd1 vccd1 vccd1 _10384_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_93_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11471_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07164_ _10023_/A0 _10343_/Q _07172_/S vssd1 vssd1 vccd1 vccd1 _07165_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11270_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06115_ _06105_/X _06106_/X _06109_/X _06114_/X vssd1 vssd1 vccd1 vccd1 _06115_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07095_ _08902_/B _07095_/B vssd1 vssd1 vccd1 vccd1 _07095_/X sky130_fd_sc_hd__or2_4
XFILLER_105_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06046_ _10701_/Q _06807_/A2 _06805_/B1 _10534_/Q _06045_/X vssd1 vssd1 vccd1 vccd1
+ _06046_/X sky130_fd_sc_hd__o221a_2
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout213 _07959_/S vssd1 vssd1 vccd1 vccd1 _07956_/S sky130_fd_sc_hd__clkbuf_4
Xfanout224 _07223_/Y vssd1 vssd1 vccd1 vccd1 _07233_/S sky130_fd_sc_hd__buf_12
Xfanout235 _10119_/X vssd1 vssd1 vccd1 vccd1 _10135_/S sky130_fd_sc_hd__buf_6
XFILLER_101_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout246 _08946_/B vssd1 vssd1 vccd1 vccd1 _08942_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09805_ _10527_/Q _09565_/A _09950_/B1 _10287_/Q vssd1 vssd1 vccd1 vccd1 _09805_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout257 _08594_/X vssd1 vssd1 vccd1 vccd1 _08621_/S sky130_fd_sc_hd__buf_6
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout268 _08272_/S vssd1 vssd1 vccd1 vccd1 _08276_/S sky130_fd_sc_hd__buf_6
XFILLER_86_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07997_ _09395_/A0 _10823_/Q _08011_/S vssd1 vssd1 vccd1 vccd1 _07998_/B sky130_fd_sc_hd__mux2_1
XFILLER_75_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout279 _07994_/X vssd1 vssd1 vccd1 vccd1 _08015_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09736_ _10340_/Q _09875_/A2 _09872_/A2 _10353_/Q _09735_/X vssd1 vssd1 vccd1 vccd1
+ _09739_/C sky130_fd_sc_hd__a221o_1
X_06948_ _09538_/A _06947_/X _06969_/S vssd1 vssd1 vccd1 vccd1 _06948_/X sky130_fd_sc_hd__mux2_4
XFILLER_86_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09667_ _11632_/Q _09434_/B _09666_/X _09678_/A vssd1 vssd1 vccd1 vccd1 _11632_/D
+ sky130_fd_sc_hd__o211a_1
X_06879_ _06874_/X _06875_/X _06878_/X _06873_/X vssd1 vssd1 vccd1 vccd1 _06879_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _08618_/A _08618_/B vssd1 vssd1 vccd1 vccd1 _11163_/D sky130_fd_sc_hd__or2_1
XFILLER_15_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09820_/A _09820_/B _09564_/A vssd1 vssd1 vccd1 vccd1 _09823_/B sky130_fd_sc_hd__a21oi_4
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08549_ _11125_/Q _08558_/S _07355_/S _07090_/A vssd1 vssd1 vccd1 vccd1 _11125_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11560_ _11810_/CLK _11560_/D vssd1 vssd1 vccd1 vccd1 _11560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10511_ _11698_/CLK _10511_/D vssd1 vssd1 vccd1 vccd1 _10511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11491_ _11495_/CLK _11491_/D vssd1 vssd1 vccd1 vccd1 _11491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10442_ _11268_/CLK _10442_/D vssd1 vssd1 vccd1 vccd1 _10442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10373_ _11706_/CLK _10373_/D vssd1 vssd1 vccd1 vccd1 _10373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout780 _09249_/A vssd1 vssd1 vccd1 vccd1 _06538_/B1 sky130_fd_sc_hd__buf_4
Xfanout791 _06737_/B1 vssd1 vssd1 vccd1 vccd1 _06717_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _05412_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _09270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_173 _07599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_184 _07070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _07021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11758_/CLK _11758_/D vssd1 vssd1 vccd1 vccd1 _11758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10709_ _11457_/CLK _10709_/D vssd1 vssd1 vccd1 vccd1 _10709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11689_ _11765_/CLK _11689_/D vssd1 vssd1 vccd1 vccd1 _11689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07920_ _07920_/A _07920_/B vssd1 vssd1 vccd1 vccd1 _10777_/D sky130_fd_sc_hd__or2_1
XFILLER_151_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07851_ _07100_/X _10744_/Q _07852_/S vssd1 vssd1 vccd1 vccd1 _10744_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_140_wb_clk_i clkbuf_4_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11177_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_151_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06802_ _11719_/Q _06857_/B1 _06801_/X _06849_/C1 vssd1 vssd1 vccd1 vccd1 _06802_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput2 io_in[6] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
X_07782_ _08684_/A _07782_/B vssd1 vssd1 vccd1 vccd1 _10698_/D sky130_fd_sc_hd__or2_1
XFILLER_49_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09521_ _09492_/B _09489_/B _09489_/C _11617_/Q vssd1 vssd1 vccd1 vccd1 _09523_/B
+ sky130_fd_sc_hd__a31o_1
X_06733_ _06728_/X _06729_/X _06730_/X _06873_/D1 vssd1 vssd1 vccd1 vccd1 _06733_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09452_ _09475_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09452_/Y sky130_fd_sc_hd__nand2_1
X_06664_ _06535_/A _06663_/X _06662_/X _06664_/C1 vssd1 vssd1 vccd1 vccd1 _06664_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ _08875_/A _08403_/B vssd1 vssd1 vccd1 vccd1 _11042_/D sky130_fd_sc_hd__or2_1
X_05615_ _05615_/A _05615_/B vssd1 vssd1 vccd1 vccd1 _05615_/Y sky130_fd_sc_hd__nor2_8
XFILLER_40_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09383_ _10183_/A0 _11550_/Q _09390_/S vssd1 vssd1 vccd1 vccd1 _11550_/D sky130_fd_sc_hd__mux2_1
X_06595_ _11179_/Q _08647_/B _06591_/X _06594_/X vssd1 vssd1 vccd1 vccd1 _06601_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_40_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08334_ _11009_/Q _08322_/Y _08325_/Y _07333_/X vssd1 vssd1 vccd1 vccd1 _11009_/D
+ sky130_fd_sc_hd__a22o_1
X_05546_ _05618_/A1 _11491_/Q _11488_/Q _05606_/B2 _05544_/X vssd1 vssd1 vccd1 vccd1
+ _05549_/A sky130_fd_sc_hd__a221o_4
XFILLER_137_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08265_ _08781_/A _08265_/B vssd1 vssd1 vccd1 vccd1 _10964_/D sky130_fd_sc_hd__or2_1
X_05477_ _10222_/Q input42/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05477_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07216_ _07034_/A _07204_/B _07771_/B1 _10373_/Q vssd1 vssd1 vccd1 vccd1 _10373_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08196_ _08196_/A _08196_/B vssd1 vssd1 vccd1 vccd1 _10933_/D sky130_fd_sc_hd__or2_1
XFILLER_118_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07147_ _07147_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _07451_/B sky130_fd_sc_hd__and2_4
XFILLER_69_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07078_ _10298_/Q _07078_/B vssd1 vssd1 vccd1 vccd1 _07078_/X sky130_fd_sc_hd__or2_1
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06029_ _11670_/Q _09965_/A _08311_/A _10995_/Q vssd1 vssd1 vccd1 vccd1 _06029_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1008 _10106_/A1 vssd1 vssd1 vccd1 vccd1 _10190_/A0 sky130_fd_sc_hd__buf_6
XFILLER_47_1374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1019 _10177_/A1 vssd1 vssd1 vccd1 vccd1 _09995_/A1 sky130_fd_sc_hd__buf_6
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09719_ _11438_/Q _09876_/A2 _09881_/B1 _10400_/Q vssd1 vssd1 vccd1 vccd1 _09719_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10991_ _11756_/CLK _10991_/D vssd1 vssd1 vccd1 vccd1 _10991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11812_/CLK _11612_/D vssd1 vssd1 vccd1 vccd1 _11612_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11543_ _11800_/CLK _11543_/D vssd1 vssd1 vccd1 vccd1 _11543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11474_ _11474_/CLK _11474_/D vssd1 vssd1 vccd1 vccd1 _11474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10425_ _11233_/CLK _10425_/D vssd1 vssd1 vccd1 vccd1 _10425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10356_ _10727_/CLK _10356_/D vssd1 vssd1 vccd1 vccd1 _10356_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_11__f_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_99_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_140_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10287_ _10812_/CLK _10287_/D vssd1 vssd1 vccd1 vccd1 _10287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05400_ _05400_/A _05400_/B _05400_/C _05400_/D vssd1 vssd1 vccd1 vccd1 _05401_/B
+ sky130_fd_sc_hd__or4_4
X_06380_ _11112_/Q _06737_/A2 _06376_/X _06379_/X vssd1 vssd1 vccd1 vccd1 _06380_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05331_ _10850_/Q _10849_/Q _05397_/S vssd1 vssd1 vccd1 vccd1 _05334_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08050_ _08050_/A _08050_/B vssd1 vssd1 vccd1 vccd1 _10851_/D sky130_fd_sc_hd__or2_1
X_05262_ _10740_/Q _10445_/Q _05397_/S vssd1 vssd1 vccd1 vccd1 _05264_/C sky130_fd_sc_hd__mux2_1
XFILLER_128_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07001_ _07205_/A _07483_/S vssd1 vssd1 vccd1 vccd1 _07044_/S sky130_fd_sc_hd__nand2_4
X_05193_ _11064_/Q _11063_/Q _06945_/B vssd1 vssd1 vccd1 vccd1 _05203_/B sky130_fd_sc_hd__mux2_1
XFILLER_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08952_ _09540_/A _08958_/A vssd1 vssd1 vccd1 vccd1 _08952_/Y sky130_fd_sc_hd__nand2_1
X_07903_ _07904_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _09208_/B sky130_fd_sc_hd__nor2_4
X_08883_ _08883_/A1 _08890_/S _08882_/X _08943_/C1 vssd1 vssd1 vccd1 vccd1 _11298_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07834_ _07025_/A _07839_/A2 _07959_/S _10729_/Q vssd1 vssd1 vccd1 vccd1 _10729_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07765_ _10685_/Q _07229_/X _07773_/S vssd1 vssd1 vccd1 vccd1 _10685_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09504_ _09522_/B _09504_/B vssd1 vssd1 vccd1 vccd1 _09504_/Y sky130_fd_sc_hd__nand2_1
X_06716_ _11121_/Q _06716_/A2 _06716_/B1 _11257_/Q vssd1 vssd1 vccd1 vccd1 _06716_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07696_ _08303_/A _08591_/B vssd1 vssd1 vccd1 vccd1 _07696_/Y sky130_fd_sc_hd__nor2_2
XFILLER_112_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09435_ _11588_/Q _11647_/Q _09440_/S vssd1 vssd1 vccd1 vccd1 _11588_/D sky130_fd_sc_hd__mux2_1
X_06647_ _10709_/Q _09059_/A _09109_/A _10544_/Q _06646_/X vssd1 vssd1 vccd1 vccd1
+ _06647_/X sky130_fd_sc_hd__a221o_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09366_ _11541_/Q _09376_/B vssd1 vssd1 vccd1 vccd1 _09366_/X sky130_fd_sc_hd__or2_1
X_06578_ _06855_/B _06577_/X _06576_/X _05730_/Y vssd1 vssd1 vccd1 vccd1 _06578_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08317_ _10114_/A0 _10996_/Q _08321_/S vssd1 vssd1 vccd1 vccd1 _10996_/D sky130_fd_sc_hd__mux2_1
X_05529_ _05631_/A2 _11507_/Q _11503_/Q _05631_/B1 _05527_/X vssd1 vssd1 vccd1 vccd1
+ _05529_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09297_ _10162_/A1 _09293_/X _09296_/X _10177_/C1 vssd1 vssd1 vccd1 vccd1 _11499_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_40 wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_62 input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_73 _05716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08248_ _10956_/Q _08284_/B vssd1 vssd1 vccd1 vccd1 _08248_/X sky130_fd_sc_hd__or2_1
XFILLER_138_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_84 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_95 _09573_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08179_ _10132_/A0 _10921_/Q _08181_/S vssd1 vssd1 vccd1 vccd1 _10921_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10210_ _11809_/CLK _10210_/D vssd1 vssd1 vccd1 vccd1 _10210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11190_ _11325_/CLK _11190_/D vssd1 vssd1 vccd1 vccd1 _11190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10141_ _11783_/Q _10137_/X _10140_/X vssd1 vssd1 vccd1 vccd1 _11783_/D sky130_fd_sc_hd__a21o_1
Xoutput180 _05477_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_4
XFILLER_47_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput191 _05478_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_4
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10072_ _10072_/A _10108_/B _10119_/C vssd1 vssd1 vccd1 vccd1 _10082_/S sky130_fd_sc_hd__or3_4
XFILLER_88_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10974_ _11572_/CLK _10974_/D vssd1 vssd1 vccd1 vccd1 _10974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11526_ _11685_/CLK _11526_/D vssd1 vssd1 vccd1 vccd1 _11526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11457_ _11457_/CLK _11457_/D vssd1 vssd1 vccd1 vccd1 _11457_/Q sky130_fd_sc_hd__dfxtp_1
X_10408_ _11470_/CLK _10408_/D vssd1 vssd1 vccd1 vccd1 _10408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11388_ _11428_/CLK _11388_/D vssd1 vssd1 vccd1 vccd1 _11388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _11471_/CLK _10339_/D vssd1 vssd1 vccd1 vccd1 _10339_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05880_ _10646_/Q _06629_/A2 _05876_/X _05879_/X vssd1 vssd1 vccd1 vccd1 _05880_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07550_ _08536_/A _07550_/B vssd1 vssd1 vccd1 vccd1 _10558_/D sky130_fd_sc_hd__or2_1
XFILLER_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06501_ _11067_/Q _06538_/A2 _06538_/B1 _11185_/Q vssd1 vssd1 vccd1 vccd1 _06501_/X
+ sky130_fd_sc_hd__o22a_1
X_07481_ _07141_/A _10519_/Q _07483_/S vssd1 vssd1 vccd1 vccd1 _07482_/B sky130_fd_sc_hd__mux2_1
X_09220_ _07187_/B _09208_/B _09205_/Y _11459_/Q _09192_/A vssd1 vssd1 vccd1 vccd1
+ _11459_/D sky130_fd_sc_hd__a221o_1
XFILLER_50_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06432_ _10403_/Q _06645_/A2 _06648_/A2 _10806_/Q vssd1 vssd1 vccd1 vccd1 _06432_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09151_ _10178_/A1 _09149_/B _10166_/B1 vssd1 vssd1 vccd1 vccd1 _09151_/X sky130_fd_sc_hd__a21o_1
X_06363_ _11487_/Q _06363_/A2 _06359_/X _06362_/X vssd1 vssd1 vccd1 vccd1 _06364_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08102_ _10875_/Q _07007_/A _08102_/S vssd1 vssd1 vccd1 vccd1 _08103_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05314_ _10609_/Q _10883_/Q _05385_/S vssd1 vssd1 vccd1 vccd1 _05318_/A sky130_fd_sc_hd__mux2_1
X_09082_ _09082_/A _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09082_/X sky130_fd_sc_hd__or3_4
X_06294_ _11496_/Q _09271_/A _06290_/X _06293_/X vssd1 vssd1 vccd1 vccd1 _06294_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_135_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08033_ _10841_/Q _08037_/B vssd1 vssd1 vccd1 vccd1 _08033_/X sky130_fd_sc_hd__or2_1
X_05245_ _10789_/Q _10863_/Q _08956_/B vssd1 vssd1 vccd1 vccd1 _05247_/C sky130_fd_sc_hd__mux2_1
Xinput60 wb_rom_val[26] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_4
Xinput71 wb_rom_val[7] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__buf_2
Xinput82 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_2
Xinput93 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__buf_2
X_05176_ _05176_/A _05176_/B _05176_/C _05176_/D vssd1 vssd1 vccd1 vccd1 _05179_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_104_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09984_ _11679_/Q _09994_/B vssd1 vssd1 vccd1 vccd1 _09984_/X sky130_fd_sc_hd__or2_1
XFILLER_44_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08935_ _08935_/A1 _08940_/S _08934_/X _08943_/C1 vssd1 vssd1 vccd1 vccd1 _11326_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08866_ _08919_/A1 _11290_/Q _08874_/S vssd1 vssd1 vccd1 vccd1 _08867_/B sky130_fd_sc_hd__mux2_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07817_ _07076_/A _10716_/Q _07817_/S vssd1 vssd1 vccd1 vccd1 _07818_/B sky130_fd_sc_hd__mux2_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08797_ _08853_/A1 _08792_/S _08796_/X _08937_/C1 vssd1 vssd1 vccd1 vccd1 _11254_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07748_ _10675_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07748_/X sky130_fd_sc_hd__or2_1
XFILLER_25_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07679_ _10635_/Q _07674_/X _07675_/Y _07090_/X vssd1 vssd1 vccd1 vccd1 _10635_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09418_ _11648_/Q _11577_/Q _09426_/S vssd1 vssd1 vccd1 vccd1 _11577_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ _10725_/CLK _10690_/D vssd1 vssd1 vccd1 vccd1 _10690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09349_ _10110_/A0 _11529_/Q _09357_/S vssd1 vssd1 vccd1 vccd1 _11529_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11311_ _11312_/CLK _11311_/D vssd1 vssd1 vccd1 vccd1 _11311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11242_ _11330_/CLK _11242_/D vssd1 vssd1 vccd1 vccd1 _11242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11173_ _11269_/CLK _11173_/D vssd1 vssd1 vccd1 vccd1 _11173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10124_ _07092_/A _11770_/Q _10135_/S vssd1 vssd1 vccd1 vccd1 _11770_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10055_ _11719_/Q _07076_/A _10057_/S vssd1 vssd1 vccd1 vccd1 _10056_/B sky130_fd_sc_hd__mux2_1
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10957_ _11683_/CLK _10957_/D vssd1 vssd1 vccd1 vccd1 _10957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10888_ _11269_/CLK _10888_/D vssd1 vssd1 vccd1 vccd1 _10888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11509_ _11735_/CLK _11509_/D vssd1 vssd1 vccd1 vccd1 _11509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout609 _06228_/A2 vssd1 vssd1 vccd1 vccd1 _06415_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06981_ _10258_/Q _06995_/B vssd1 vssd1 vccd1 vccd1 _06981_/X sky130_fd_sc_hd__or2_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05932_ _11125_/Q _06635_/A2 _05931_/X _06550_/C1 vssd1 vssd1 vccd1 vccd1 _05932_/X
+ sky130_fd_sc_hd__o211a_1
X_08720_ _11216_/Q _08726_/S _07852_/S _07098_/B vssd1 vssd1 vccd1 vccd1 _11216_/D
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11809_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08651_ _11181_/Q _08655_/B _08750_/B vssd1 vssd1 vccd1 vccd1 _08651_/X sky130_fd_sc_hd__or3_1
X_05863_ _10456_/Q _06643_/A2 _06640_/B1 _11136_/Q _05860_/X vssd1 vssd1 vccd1 vccd1
+ _05864_/C sky130_fd_sc_hd__o221a_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07602_ _10582_/Q _07598_/Y _07599_/Y _08441_/B2 vssd1 vssd1 vccd1 vccd1 _10582_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_54_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08582_ _09395_/A0 _08589_/S _08581_/X _08588_/C1 vssd1 vssd1 vccd1 vccd1 _11146_/D
+ sky130_fd_sc_hd__o211a_1
X_05794_ _11069_/Q _06731_/B1 _07111_/A _11766_/Q vssd1 vssd1 vccd1 vccd1 _05794_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07533_ _07076_/A _10551_/Q _07533_/S vssd1 vssd1 vccd1 vccd1 _07534_/B sky130_fd_sc_hd__mux2_1
XFILLER_74_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07464_ _07476_/A _07464_/B vssd1 vssd1 vccd1 vccd1 _10509_/D sky130_fd_sc_hd__or2_1
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09203_ _11449_/Q _09190_/Y _09193_/Y _07040_/X vssd1 vssd1 vccd1 vccd1 _11449_/D
+ sky130_fd_sc_hd__a22o_1
X_06415_ _10828_/Q _06415_/A2 _06628_/B1 _11273_/Q vssd1 vssd1 vccd1 vccd1 _06415_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07395_ _07048_/A _10474_/Q _07429_/S vssd1 vssd1 vccd1 vccd1 _07396_/B sky130_fd_sc_hd__mux2_1
X_09134_ _10161_/A1 _09132_/X _09133_/X _09168_/C1 vssd1 vssd1 vccd1 vccd1 _11412_/D
+ sky130_fd_sc_hd__o211a_1
X_06346_ _11765_/Q _10108_/A _06344_/X _06345_/X vssd1 vssd1 vccd1 vccd1 _06346_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09065_ _11381_/Q _09077_/B vssd1 vssd1 vccd1 vccd1 _09065_/X sky130_fd_sc_hd__or2_1
XFILLER_50_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06277_ _06450_/A _10229_/Q _08970_/S _06276_/X vssd1 vssd1 vccd1 vccd1 _10229_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08016_ _08833_/A _08016_/B vssd1 vssd1 vccd1 vccd1 _10832_/D sky130_fd_sc_hd__or2_1
X_05228_ _05419_/S _11010_/Q vssd1 vssd1 vccd1 vccd1 _05228_/X sky130_fd_sc_hd__and2b_1
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05159_ _11080_/Q _10600_/Q _05399_/S vssd1 vssd1 vccd1 vccd1 _05162_/B sky130_fd_sc_hd__mux2_1
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09967_ _10110_/A0 _11667_/Q _09975_/S vssd1 vssd1 vccd1 vccd1 _11667_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08918_ _11318_/Q _08946_/B vssd1 vssd1 vccd1 vccd1 _08918_/X sky130_fd_sc_hd__or2_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _11702_/Q _09571_/B _09566_/A _11696_/Q _09897_/X vssd1 vssd1 vccd1 vccd1
+ _09899_/D sky130_fd_sc_hd__a221o_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08849_ _08935_/A1 _08850_/S _08848_/X _07011_/B vssd1 vssd1 vccd1 vccd1 _11282_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ _10812_/CLK _10811_/D vssd1 vssd1 vccd1 vccd1 _10811_/Q sky130_fd_sc_hd__dfxtp_1
X_11791_ _11791_/CLK _11791_/D vssd1 vssd1 vccd1 vccd1 _11791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10742_ _11262_/CLK _10742_/D vssd1 vssd1 vccd1 vccd1 _10742_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10673_ _10782_/CLK _10673_/D vssd1 vssd1 vccd1 vccd1 _10673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11225_ _11651_/CLK _11225_/D vssd1 vssd1 vccd1 vccd1 _11225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11156_ _11251_/CLK _11156_/D vssd1 vssd1 vccd1 vccd1 _11156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10107_ _11755_/Q _10087_/X _10106_/X vssd1 vssd1 vccd1 vccd1 _11755_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11087_ _11607_/CLK _11087_/D vssd1 vssd1 vccd1 vccd1 _11087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10038_ _11709_/Q _10134_/A0 _10051_/S vssd1 vssd1 vccd1 vccd1 _10039_/B sky130_fd_sc_hd__mux2_1
XFILLER_36_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06200_ _06190_/X _06191_/X _06194_/X _06199_/X vssd1 vssd1 vccd1 vccd1 _06200_/X
+ sky130_fd_sc_hd__a31o_4
X_07180_ _07034_/A _10351_/Q _09240_/S vssd1 vssd1 vccd1 vccd1 _07181_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06131_ _06127_/X _06130_/X _07083_/A _06125_/X vssd1 vssd1 vccd1 vccd1 _06131_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_121_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06062_ _10464_/Q _06371_/A2 _07827_/A2 _10979_/Q vssd1 vssd1 vccd1 vccd1 _06062_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout406 _05390_/Y vssd1 vssd1 vccd1 vccd1 _09947_/B1 sky130_fd_sc_hd__buf_6
Xfanout417 _05335_/Y vssd1 vssd1 vccd1 vccd1 _09882_/B1 sky130_fd_sc_hd__buf_4
XFILLER_59_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09821_ _09515_/B _09820_/X _09824_/S vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout428 _09572_/A vssd1 vssd1 vccd1 vccd1 _09953_/B1 sky130_fd_sc_hd__buf_6
XFILLER_87_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout439 _05214_/Y vssd1 vssd1 vccd1 vccd1 _09875_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09752_ _10503_/Q _09871_/A2 _09886_/B1 _10552_/Q _09751_/X vssd1 vssd1 vccd1 vccd1
+ _09757_/B sky130_fd_sc_hd__a221o_1
X_06964_ _05474_/A _06962_/X _06963_/X _06950_/A vssd1 vssd1 vccd1 vccd1 _06964_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08703_ _11206_/Q _08705_/B vssd1 vssd1 vccd1 vccd1 _08703_/X sky130_fd_sc_hd__or2_1
X_05915_ _10699_/Q _07778_/A _06805_/B1 _10497_/Q _05914_/X vssd1 vssd1 vccd1 vccd1
+ _05915_/X sky130_fd_sc_hd__o221a_1
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09683_ _11639_/Q _09692_/B vssd1 vssd1 vccd1 vccd1 _09683_/X sky130_fd_sc_hd__or2_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06895_ _06901_/A _08243_/C _08243_/D vssd1 vssd1 vccd1 vccd1 _10180_/B sky130_fd_sc_hd__or3_4
XFILLER_67_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05846_ _10281_/Q _07046_/A _06238_/A2 _10475_/Q _05845_/X vssd1 vssd1 vccd1 vccd1
+ _05846_/X sky130_fd_sc_hd__o221a_1
X_08634_ _07070_/A _08621_/S _08633_/X _07003_/B vssd1 vssd1 vccd1 vccd1 _11171_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05777_ _10280_/Q _07046_/A _07190_/A _10474_/Q _05776_/X vssd1 vssd1 vccd1 vccd1
+ _05777_/X sky130_fd_sc_hd__o221a_1
X_08565_ _11136_/Q _08577_/S _08563_/Y _07005_/A vssd1 vssd1 vccd1 vccd1 _11136_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07516_ _07818_/A _07516_/B vssd1 vssd1 vccd1 vccd1 _10542_/D sky130_fd_sc_hd__or2_1
XFILLER_126_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08496_ _08664_/A _08496_/B vssd1 vssd1 vccd1 vccd1 _11098_/D sky130_fd_sc_hd__or2_1
XFILLER_74_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07447_ _09214_/A _07533_/S _07442_/Y _10499_/Q _09193_/A vssd1 vssd1 vccd1 vccd1
+ _10499_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07378_ _08745_/A _07378_/B vssd1 vssd1 vccd1 vccd1 _10463_/D sky130_fd_sc_hd__or2_1
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09117_ _10166_/A1 _09127_/B _09129_/B1 vssd1 vssd1 vccd1 vccd1 _09117_/X sky130_fd_sc_hd__a21o_1
X_06329_ _10468_/Q _06642_/A2 _08469_/B _11081_/Q vssd1 vssd1 vccd1 vccd1 _06329_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09048_ _09280_/A1 _09038_/X _09047_/X _09048_/C1 vssd1 vssd1 vccd1 vccd1 _11373_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _11235_/CLK _11010_/D vssd1 vssd1 vccd1 vccd1 _11010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout940 _09237_/A0 vssd1 vssd1 vccd1 vccd1 _07028_/A sky130_fd_sc_hd__buf_6
Xfanout951 fanout958/X vssd1 vssd1 vccd1 vccd1 _08818_/A1 sky130_fd_sc_hd__buf_8
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout962 input92/X vssd1 vssd1 vccd1 vccd1 _08935_/A1 sky130_fd_sc_hd__buf_6
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout973 input89/X vssd1 vssd1 vccd1 vccd1 _08969_/A1 sky130_fd_sc_hd__clkbuf_8
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout984 input85/X vssd1 vssd1 vccd1 vccd1 _11872_/A sky130_fd_sc_hd__buf_12
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 _06357_/C1 vssd1 vssd1 vccd1 vccd1 _07298_/B sky130_fd_sc_hd__clkbuf_16
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1086 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1086/HI io_oeb[16] sky130_fd_sc_hd__conb_1
XFILLER_57_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1097 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1097/HI io_oeb[27] sky130_fd_sc_hd__conb_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11774_ _11779_/CLK _11774_/D vssd1 vssd1 vccd1 vccd1 _11774_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _10725_/CLK _10725_/D vssd1 vssd1 vccd1 vccd1 _10725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10656_ _11442_/CLK _10656_/D vssd1 vssd1 vccd1 vccd1 _10656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10587_ _11243_/CLK _10587_/D vssd1 vssd1 vccd1 vccd1 _10587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ _11319_/CLK _11208_/D vssd1 vssd1 vccd1 vccd1 _11208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11139_ _11651_/CLK _11139_/D vssd1 vssd1 vccd1 vccd1 _11139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05700_ _11111_/Q _05549_/Y _05555_/Y _11114_/Q _05699_/X vssd1 vssd1 vccd1 vccd1
+ _05703_/B sky130_fd_sc_hd__a221o_1
X_06680_ _11119_/Q _06737_/A2 _06677_/X _06679_/X vssd1 vssd1 vccd1 vccd1 _06680_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05631_ _11791_/Q _05631_/A2 _05631_/B1 _11787_/Q _05629_/X vssd1 vssd1 vccd1 vccd1
+ _05631_/X sky130_fd_sc_hd__a221o_1
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08350_ _11018_/Q _08362_/B vssd1 vssd1 vccd1 vccd1 _08350_/X sky130_fd_sc_hd__or2_1
X_05562_ _11799_/Q _05616_/A1 _05077_/A _11796_/Q vssd1 vssd1 vccd1 vccd1 _05562_/X
+ sky130_fd_sc_hd__a22o_1
X_07301_ _08322_/A _08762_/B vssd1 vssd1 vccd1 vccd1 _07301_/Y sky130_fd_sc_hd__nor2_2
XFILLER_32_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08281_ _09237_/A0 _08272_/S _08280_/X _07003_/B vssd1 vssd1 vccd1 vccd1 _10972_/D
+ sky130_fd_sc_hd__o211a_1
X_05493_ _10238_/Q input49/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05493_/X sky130_fd_sc_hd__mux2_1
X_07232_ _08655_/B _07232_/B vssd1 vssd1 vccd1 vccd1 _07232_/X sky130_fd_sc_hd__or2_4
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07163_ _07920_/A _07163_/B vssd1 vssd1 vccd1 vccd1 _10342_/D sky130_fd_sc_hd__or2_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06114_ _10771_/Q _06862_/A2 _06110_/X _06113_/X vssd1 vssd1 vccd1 vccd1 _06114_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_106_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07094_ _10302_/Q _07093_/X _07109_/S vssd1 vssd1 vccd1 vccd1 _10302_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06045_ _10398_/Q _06804_/B _07540_/A _10558_/Q vssd1 vssd1 vccd1 vccd1 _06045_/X
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_62_wb_clk_i clkbuf_leaf_69_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11527_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout214 _07959_/S vssd1 vssd1 vccd1 vccd1 _07961_/S sky130_fd_sc_hd__buf_6
Xfanout225 _07205_/Y vssd1 vssd1 vccd1 vccd1 _07773_/S sky130_fd_sc_hd__buf_6
Xfanout236 _10119_/X vssd1 vssd1 vccd1 vccd1 _10134_/S sky130_fd_sc_hd__buf_4
X_09804_ _10295_/Q _09570_/A _09570_/B _10292_/Q vssd1 vssd1 vccd1 vccd1 _09804_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout247 _08906_/Y vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__buf_4
Xfanout258 _08594_/X vssd1 vssd1 vccd1 vccd1 _08623_/S sky130_fd_sc_hd__buf_6
Xfanout269 _08245_/X vssd1 vssd1 vccd1 vccd1 _08272_/S sky130_fd_sc_hd__buf_8
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07996_ _07007_/A _08011_/S _07995_/X _08831_/C1 vssd1 vssd1 vccd1 vccd1 _10822_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09735_ _10343_/Q _09877_/A2 _09886_/B1 _11473_/Q vssd1 vssd1 vccd1 vccd1 _09735_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06947_ _11605_/Q _09538_/C _06944_/A _08955_/A vssd1 vssd1 vccd1 vccd1 _06947_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09666_ _11634_/Q _09540_/A _09692_/B _11629_/Q vssd1 vssd1 vccd1 vccd1 _09666_/X
+ sky130_fd_sc_hd__a211o_1
X_06878_ _11450_/Q _07777_/A _06877_/X _06878_/C1 vssd1 vssd1 vccd1 vccd1 _06878_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08617_ _08789_/A1 _11163_/Q _08621_/S vssd1 vssd1 vccd1 vccd1 _08618_/B sky130_fd_sc_hd__mux2_1
X_05829_ _11390_/Q _09082_/A _06716_/B1 _11403_/Q vssd1 vssd1 vccd1 vccd1 _05829_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09597_ _11643_/Q _09596_/B _09594_/X vssd1 vssd1 vccd1 vccd1 _09820_/B sky130_fd_sc_hd__a21o_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08548_ _11124_/Q _08558_/S _07357_/S _07005_/A vssd1 vssd1 vccd1 vccd1 _11124_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08479_ _11090_/Q _08503_/B vssd1 vssd1 vccd1 vccd1 _08479_/X sky130_fd_sc_hd__or2_1
XFILLER_126_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10510_ _11702_/CLK _10510_/D vssd1 vssd1 vccd1 vccd1 _10510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11490_ _11497_/CLK _11490_/D vssd1 vssd1 vccd1 vccd1 _11490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10441_ _11268_/CLK _10441_/D vssd1 vssd1 vccd1 vccd1 _10441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10372_ _11745_/CLK _10372_/D vssd1 vssd1 vccd1 vccd1 _10372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_10__f_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout770 _10119_/A vssd1 vssd1 vccd1 vccd1 _06639_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_77_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout781 fanout782/X vssd1 vssd1 vccd1 vccd1 _09249_/A sky130_fd_sc_hd__clkbuf_4
Xfanout792 fanout793/X vssd1 vssd1 vccd1 vccd1 _06737_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _07018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _05434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_152 _07052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _05432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _07070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_196 _07015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _11763_/CLK _11757_/D vssd1 vssd1 vccd1 vccd1 _11757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10708_ _10782_/CLK _10708_/D vssd1 vssd1 vccd1 vccd1 _10708_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11688_ _11735_/CLK _11688_/D vssd1 vssd1 vccd1 vccd1 _11688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10639_ _10644_/CLK _10639_/D vssd1 vssd1 vccd1 vccd1 _10639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07850_ _08441_/B2 _10743_/Q _07852_/S vssd1 vssd1 vccd1 vccd1 _10743_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06801_ _10297_/Q _06106_/B _06871_/B1 _10801_/Q _06800_/X vssd1 vssd1 vccd1 vccd1
+ _06801_/X sky130_fd_sc_hd__o221a_1
XFILLER_151_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07781_ _10013_/A0 _10698_/Q _07817_/S vssd1 vssd1 vccd1 vccd1 _07782_/B sky130_fd_sc_hd__mux2_1
Xinput3 io_in[7] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09520_ _09525_/A _09486_/X _09528_/B _09519_/X _09529_/A vssd1 vssd1 vccd1 vccd1
+ _11616_/D sky130_fd_sc_hd__o311a_1
X_06732_ _10294_/Q _07046_/A _07111_/A _10328_/Q _06731_/X vssd1 vssd1 vccd1 vccd1
+ _06732_/X sky130_fd_sc_hd__o221a_2
XFILLER_37_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06663_ _06663_/A _10237_/Q vssd1 vssd1 vccd1 vccd1 _06663_/X sky130_fd_sc_hd__and2_1
X_09451_ input32/X _09442_/X _09450_/X vssd1 vssd1 vccd1 vccd1 _09452_/B sky130_fd_sc_hd__o21ai_1
XFILLER_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05614_ _11627_/Q _11395_/Q _11390_/Q _05620_/B2 _05613_/X vssd1 vssd1 vccd1 vccd1
+ _05615_/B sky130_fd_sc_hd__a221o_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08402_ _09101_/A1 _11042_/Q _08404_/S vssd1 vssd1 vccd1 vccd1 _08403_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09382_ _10110_/A0 _11549_/Q _09390_/S vssd1 vssd1 vccd1 vccd1 _11549_/D sky130_fd_sc_hd__mux2_1
X_06594_ _10600_/Q _06636_/A2 _06593_/X _11869_/A vssd1 vssd1 vccd1 vccd1 _06594_/X
+ sky130_fd_sc_hd__o211a_1
X_05545_ _09552_/A1 _11496_/Q _11490_/Q _05078_/A vssd1 vssd1 vccd1 vccd1 _05545_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08333_ _11008_/Q _08323_/Y _08324_/Y _07318_/X vssd1 vssd1 vccd1 vccd1 _11008_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08264_ _09101_/A1 _10964_/Q _08272_/S vssd1 vssd1 vccd1 vccd1 _08265_/B sky130_fd_sc_hd__mux2_1
X_05476_ input77/X input78/X vssd1 vssd1 vccd1 vccd1 _05508_/S sky130_fd_sc_hd__nor2_8
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07215_ _10047_/A1 _07205_/B _07772_/S _10372_/Q vssd1 vssd1 vccd1 vccd1 _10372_/D
+ sky130_fd_sc_hd__o22a_1
X_08195_ _10933_/Q _08818_/A1 _08197_/S vssd1 vssd1 vccd1 vccd1 _08196_/B sky130_fd_sc_hd__mux2_1
XFILLER_134_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07146_ _07036_/A _07111_/X _07145_/X _07141_/B vssd1 vssd1 vccd1 vccd1 _10334_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07077_ _10297_/Q _07045_/Y _07496_/S _07187_/B vssd1 vssd1 vccd1 vccd1 _10297_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06028_ _06024_/X _06027_/X _07297_/A _06022_/X vssd1 vssd1 vccd1 vccd1 _06028_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1009 _07057_/A vssd1 vssd1 vccd1 vccd1 _10106_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_87_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ _10813_/Q _07977_/S _07363_/S _07617_/B vssd1 vssd1 vccd1 vccd1 _10813_/D
+ sky130_fd_sc_hd__o22a_1
X_09718_ _10413_/Q _09872_/A2 _09884_/A2 _11435_/Q _09717_/X vssd1 vssd1 vccd1 vccd1
+ _09721_/C sky130_fd_sc_hd__a221o_1
XFILLER_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ _11633_/CLK _10990_/D vssd1 vssd1 vccd1 vccd1 _10990_/Q sky130_fd_sc_hd__dfxtp_1
X_09649_ _10333_/Q _09572_/C _09573_/D _10316_/Q _09648_/X vssd1 vssd1 vccd1 vccd1
+ _09650_/D sky130_fd_sc_hd__a221o_1
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11622_/CLK _11611_/D vssd1 vssd1 vccd1 vccd1 _11611_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_93_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ _11801_/CLK _11542_/D vssd1 vssd1 vccd1 vccd1 _11542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11473_ _11473_/CLK _11473_/D vssd1 vssd1 vccd1 vccd1 _11473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10424_ _10644_/CLK _10424_/D vssd1 vssd1 vccd1 vccd1 _10424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10355_ _11698_/CLK _10355_/D vssd1 vssd1 vccd1 vccd1 _10355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10812_/CLK _10286_/D vssd1 vssd1 vccd1 vccd1 _10286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11809_ _11809_/CLK _11809_/D vssd1 vssd1 vccd1 vccd1 _11809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05330_ _10456_/Q _10455_/Q _05391_/S vssd1 vssd1 vccd1 vccd1 _05334_/A sky130_fd_sc_hd__mux2_1
X_05261_ _10446_/Q _10741_/Q _05399_/S vssd1 vssd1 vccd1 vccd1 _05264_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07000_ _10039_/A _07000_/B vssd1 vssd1 vccd1 vccd1 _07000_/Y sky130_fd_sc_hd__nor2_4
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05192_ _11028_/Q _11027_/Q _05416_/S vssd1 vssd1 vccd1 vccd1 _05203_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08951_ _09554_/A _11604_/Q _11603_/Q vssd1 vssd1 vccd1 vccd1 _08951_/X sky130_fd_sc_hd__or3b_4
XFILLER_29_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07902_ _07042_/A _07966_/S _07901_/X _07902_/C1 vssd1 vssd1 vccd1 vccd1 _10769_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08882_ _11298_/Q _08894_/B vssd1 vssd1 vccd1 vccd1 _08882_/X sky130_fd_sc_hd__or2_1
XFILLER_96_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07833_ _07211_/A _07820_/B _07821_/A _10728_/Q vssd1 vssd1 vccd1 vccd1 _10728_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07764_ _10684_/Q _07227_/X _07773_/S vssd1 vssd1 vccd1 vccd1 _10684_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09503_ _11611_/Q _09501_/Y _09502_/X _09529_/A vssd1 vssd1 vccd1 vccd1 _11611_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06715_ _06709_/X _06714_/X _06743_/B vssd1 vssd1 vccd1 vccd1 _06715_/Y sky130_fd_sc_hd__o21ai_2
X_07695_ _07303_/X _08589_/S _07694_/Y _10645_/Q _08427_/A vssd1 vssd1 vccd1 vccd1
+ _10645_/D sky130_fd_sc_hd__o221a_1
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09434_ _09678_/A _09434_/B vssd1 vssd1 vccd1 vccd1 _09440_/S sky130_fd_sc_hd__and2_4
X_06646_ _10779_/Q _06646_/A2 _09131_/A _10668_/Q vssd1 vssd1 vccd1 vccd1 _06646_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09365_ _11540_/Q _09359_/X _09364_/X vssd1 vssd1 vccd1 vccd1 _11540_/D sky130_fd_sc_hd__a21o_1
X_06577_ _06577_/A _10235_/Q vssd1 vssd1 vccd1 vccd1 _06577_/X sky130_fd_sc_hd__and2_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08316_ _10113_/A0 _10995_/Q _08321_/S vssd1 vssd1 vccd1 vccd1 _10995_/D sky130_fd_sc_hd__mux2_1
X_05528_ _05618_/A1 _11501_/Q _11498_/Q _05606_/B2 _05526_/X vssd1 vssd1 vccd1 vccd1
+ _05531_/A sky130_fd_sc_hd__a221o_4
X_09296_ _11499_/Q _09310_/B vssd1 vssd1 vccd1 vccd1 _09296_/X sky130_fd_sc_hd__or2_1
XANTENNA_30 _07095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 _10233_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05459_ _10760_/Q _09883_/B1 _09950_/B1 _10753_/Q vssd1 vssd1 vccd1 vccd1 _05459_/X
+ sky130_fd_sc_hd__a22o_1
X_08247_ _09111_/A1 _08276_/S _08246_/X _08919_/C1 vssd1 vssd1 vccd1 vccd1 _10955_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_74 _11611_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_85 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 _09572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08178_ _07061_/A _10920_/Q _08181_/S vssd1 vssd1 vccd1 vccd1 _10920_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07129_ _07211_/A _07111_/X _07128_/X _07141_/B vssd1 vssd1 vccd1 vccd1 _10324_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10140_ _10182_/A0 _10154_/B _10156_/B1 vssd1 vssd1 vccd1 vccd1 _10140_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput170 _11868_/X vssd1 vssd1 vccd1 vccd1 wb_rom_adrb[2] sky130_fd_sc_hd__buf_4
Xoutput181 _05487_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_4
Xoutput192 _05497_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_4
X_10071_ _10118_/A0 _11732_/Q _10071_/S vssd1 vssd1 vccd1 vccd1 _11732_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10973_ _11291_/CLK _10973_/D vssd1 vssd1 vccd1 vccd1 _10973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11525_ _11683_/CLK _11525_/D vssd1 vssd1 vccd1 vccd1 _11525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11456_ _11471_/CLK _11456_/D vssd1 vssd1 vccd1 vccd1 _11456_/Q sky130_fd_sc_hd__dfxtp_2
X_10407_ _10808_/CLK _10407_/D vssd1 vssd1 vccd1 vccd1 _10407_/Q sky130_fd_sc_hd__dfxtp_2
X_11387_ _11428_/CLK _11387_/D vssd1 vssd1 vccd1 vccd1 _11387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10338_ _10765_/CLK _10338_/D vssd1 vssd1 vccd1 vccd1 _10338_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11744_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _11661_/CLK _10269_/D vssd1 vssd1 vccd1 vccd1 _10269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06500_ _10857_/Q _06631_/A2 _06496_/X _06499_/X vssd1 vssd1 vccd1 vccd1 _06500_/X
+ sky130_fd_sc_hd__o211a_1
X_07480_ _10043_/A _07480_/B vssd1 vssd1 vccd1 vccd1 _10518_/D sky130_fd_sc_hd__or2_1
XFILLER_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06431_ _06431_/A _06431_/B _06431_/C vssd1 vssd1 vccd1 vccd1 _06431_/X sky130_fd_sc_hd__or3_4
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09150_ _09172_/A1 _09132_/X _09149_/X _10175_/C1 vssd1 vssd1 vccd1 vccd1 _11420_/D
+ sky130_fd_sc_hd__o211a_1
X_06362_ _11801_/Q _10159_/A _06361_/X _06624_/C1 vssd1 vssd1 vccd1 vccd1 _06362_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08101_ _07232_/B _08362_/B _08100_/X vssd1 vssd1 vccd1 vccd1 _10874_/D sky130_fd_sc_hd__a21o_1
X_05313_ _05313_/A _05313_/B vssd1 vssd1 vccd1 vccd1 _05313_/Y sky130_fd_sc_hd__nor2_8
X_06293_ _11377_/Q _09038_/A _06292_/X _06357_/C1 vssd1 vssd1 vccd1 vccd1 _06293_/X
+ sky130_fd_sc_hd__o211a_1
X_09081_ _09081_/A _10136_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09099_/B sky130_fd_sc_hd__and3_4
X_08032_ _08847_/A _08032_/B vssd1 vssd1 vccd1 vccd1 _10840_/D sky130_fd_sc_hd__or2_1
X_05244_ _10792_/Q _10791_/Q _06945_/B vssd1 vssd1 vccd1 vccd1 _05247_/B sky130_fd_sc_hd__mux2_1
XFILLER_135_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput50 wb_rom_val[17] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_4
Xinput61 wb_rom_val[27] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput72 wb_rom_val[8] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_2
Xinput83 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__buf_2
Xinput94 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__buf_8
X_05175_ _11222_/Q _11221_/Q _05396_/S vssd1 vssd1 vccd1 vccd1 _05176_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09983_ _11678_/Q _09977_/X _09982_/X vssd1 vssd1 vccd1 vccd1 _11678_/D sky130_fd_sc_hd__a21o_1
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08934_ _11326_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08934_/X sky130_fd_sc_hd__or2_1
XFILLER_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08865_ _09280_/A1 _08890_/S _08864_/X _09122_/C1 vssd1 vssd1 vccd1 vccd1 _11289_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07816_ _07936_/A _07816_/B vssd1 vssd1 vccd1 vccd1 _10715_/D sky130_fd_sc_hd__or2_1
XFILLER_84_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08796_ _11254_/Q _08804_/B vssd1 vssd1 vccd1 vccd1 _08796_/X sky130_fd_sc_hd__or2_1
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07747_ _07034_/A _07751_/A2 _07746_/X _09201_/A1 vssd1 vssd1 vccd1 vccd1 _10674_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07678_ _10634_/Q _07674_/X _07675_/Y _07225_/X vssd1 vssd1 vccd1 vccd1 _10634_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09417_ _11647_/Q _11576_/Q _09704_/B vssd1 vssd1 vccd1 vccd1 _11576_/D sky130_fd_sc_hd__mux2_1
X_06629_ _11151_/Q _06629_/A2 _06629_/B1 _11102_/Q _07298_/B vssd1 vssd1 vccd1 vccd1
+ _06629_/X sky130_fd_sc_hd__o221a_2
XFILLER_12_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09348_ _09999_/A0 _11528_/Q _09357_/S vssd1 vssd1 vccd1 vccd1 _11528_/D sky130_fd_sc_hd__mux2_1
XFILLER_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09279_ _10166_/A1 _09271_/X _09278_/X _09279_/C1 vssd1 vssd1 vccd1 vccd1 _11491_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _11310_/CLK _11310_/D vssd1 vssd1 vccd1 vccd1 _11310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11241_ _11683_/CLK _11241_/D vssd1 vssd1 vccd1 vccd1 _11241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11172_ _11632_/CLK _11172_/D vssd1 vssd1 vccd1 vccd1 _11172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ _07010_/A _11769_/Q _10135_/S vssd1 vssd1 vccd1 vccd1 _11769_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10054_ _10058_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _11718_/D sky130_fd_sc_hd__or2_1
XFILLER_0_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10956_ _11393_/CLK _10956_/D vssd1 vssd1 vccd1 vccd1 _10956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10887_ _10929_/CLK _10887_/D vssd1 vssd1 vccd1 vccd1 _10887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11508_ _11756_/CLK _11508_/D vssd1 vssd1 vccd1 vccd1 _11508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11439_ _11439_/CLK _11439_/D vssd1 vssd1 vccd1 vccd1 _11439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _10182_/A0 _06976_/X _06979_/X _06990_/C1 vssd1 vssd1 vccd1 vccd1 _10257_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05931_ _11209_/Q _06637_/A2 _08647_/B _10301_/Q _05930_/X vssd1 vssd1 vccd1 vccd1
+ _05931_/X sky130_fd_sc_hd__o221a_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08650_ _08650_/A _10180_/C _10119_/B vssd1 vssd1 vccd1 vccd1 _08650_/X sky130_fd_sc_hd__or3_2
X_05862_ _10608_/Q _06468_/B _06152_/B _10611_/Q _06642_/C1 vssd1 vssd1 vccd1 vccd1
+ _05864_/B sky130_fd_sc_hd__o221a_1
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07601_ _10581_/Q _07597_/Y _07600_/Y _08440_/B2 vssd1 vssd1 vccd1 vccd1 _10581_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08581_ _11146_/Q _08591_/B vssd1 vssd1 vccd1 vccd1 _08581_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_87_wb_clk_i clkbuf_leaf_88_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11663_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05793_ _11033_/Q _09060_/A _05788_/X _05792_/X vssd1 vssd1 vccd1 vccd1 _05793_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07532_ _07926_/A _07532_/B vssd1 vssd1 vccd1 vccd1 _10550_/D sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11224_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07463_ _07052_/A _10509_/Q _07477_/S vssd1 vssd1 vccd1 vccd1 _07464_/B sky130_fd_sc_hd__mux2_1
X_09202_ _11448_/Q _09190_/Y _09193_/Y _07451_/X vssd1 vssd1 vccd1 vccd1 _11448_/D
+ sky130_fd_sc_hd__a22o_1
X_06414_ _11007_/Q _06504_/B1 _06410_/X _06413_/X vssd1 vssd1 vccd1 vccd1 _06420_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07394_ _08578_/A _07394_/B vssd1 vssd1 vccd1 vccd1 _10473_/D sky130_fd_sc_hd__and2_1
XFILLER_50_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ _11412_/Q _09149_/B vssd1 vssd1 vccd1 vccd1 _09133_/X sky130_fd_sc_hd__or2_1
X_06345_ _11732_/Q _10061_/A _09347_/A _11537_/Q vssd1 vssd1 vccd1 vccd1 _06345_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09064_ _09275_/A1 _09060_/X _09063_/X _09078_/C1 vssd1 vssd1 vccd1 vccd1 _11380_/D
+ sky130_fd_sc_hd__o211a_1
X_06276_ _05728_/X _06622_/A2 _06274_/X _06275_/Y vssd1 vssd1 vccd1 vccd1 _06276_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08015_ _08818_/A1 _10832_/Q _08015_/S vssd1 vssd1 vccd1 vccd1 _08016_/B sky130_fd_sc_hd__mux2_1
X_05227_ _11006_/Q _11005_/Q _05300_/S vssd1 vssd1 vccd1 vccd1 _05237_/B sky130_fd_sc_hd__mux2_1
XFILLER_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05158_ _11076_/Q _11075_/Q _05392_/S vssd1 vssd1 vccd1 vccd1 _05162_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09966_ _09999_/A0 _11666_/Q _09975_/S vssd1 vssd1 vccd1 vccd1 _11666_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05089_ _11032_/Q vssd1 vssd1 vccd1 vccd1 _08380_/A sky130_fd_sc_hd__inv_2
XFILLER_89_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08917_ _09280_/A1 _08940_/S _08916_/X _08943_/C1 vssd1 vssd1 vccd1 vccd1 _11317_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _11711_/Q _09565_/A _09570_/B _11712_/Q vssd1 vssd1 vccd1 vccd1 _09897_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08848_ _11282_/Q _08852_/B vssd1 vssd1 vccd1 vccd1 _08848_/X sky130_fd_sc_hd__or2_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _09124_/A1 _08802_/S _08778_/X _08947_/C1 vssd1 vssd1 vccd1 vccd1 _11245_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10810_ _11308_/CLK _10810_/D vssd1 vssd1 vccd1 vccd1 _10810_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11791_/CLK _11790_/D vssd1 vssd1 vccd1 vccd1 _11790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10741_ _11780_/CLK _10741_/D vssd1 vssd1 vccd1 vccd1 _10741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10672_ _11457_/CLK _10672_/D vssd1 vssd1 vccd1 vccd1 _10672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11224_ _11224_/CLK _11224_/D vssd1 vssd1 vccd1 vccd1 _11224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11155_ _11330_/CLK _11155_/D vssd1 vssd1 vccd1 vccd1 _11155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10106_ _10106_/A1 _10104_/B _10156_/B1 vssd1 vssd1 vccd1 vccd1 _10106_/X sky130_fd_sc_hd__a21o_1
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11086_ _11651_/CLK _11086_/D vssd1 vssd1 vccd1 vccd1 _11086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10037_ _10039_/A _10037_/B vssd1 vssd1 vccd1 vccd1 _11708_/D sky130_fd_sc_hd__or2_1
XFILLER_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10939_ _10939_/CLK _10939_/D vssd1 vssd1 vccd1 vccd1 _10939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06130_ _11260_/Q _07190_/A _06128_/X _06129_/X vssd1 vssd1 vccd1 vccd1 _06130_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_134_wb_clk_i clkbuf_4_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11706_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_06061_ _10877_/Q _06513_/A2 _06636_/A2 _10925_/Q _07083_/B vssd1 vssd1 vccd1 vccd1
+ _06061_/X sky130_fd_sc_hd__o221a_4
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout407 _05390_/Y vssd1 vssd1 vccd1 vccd1 _09565_/D sky130_fd_sc_hd__clkbuf_8
X_09820_ _09820_/A _09820_/B vssd1 vssd1 vccd1 vccd1 _09820_/X sky130_fd_sc_hd__xor2_2
Xfanout418 _05324_/Y vssd1 vssd1 vccd1 vccd1 _09573_/C sky130_fd_sc_hd__buf_8
XFILLER_119_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout429 _05270_/Y vssd1 vssd1 vccd1 vccd1 _09572_/A sky130_fd_sc_hd__buf_6
XFILLER_28_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09751_ _10501_/Q _09883_/B1 _09565_/D _10546_/Q _09750_/X vssd1 vssd1 vccd1 vccd1
+ _09751_/X sky130_fd_sc_hd__a221o_1
XFILLER_100_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06963_ _09538_/B input8/X _09488_/C vssd1 vssd1 vccd1 vccd1 _06963_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08702_ _09216_/A0 _08707_/S _08701_/X _08937_/C1 vssd1 vssd1 vccd1 vccd1 _11205_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05914_ _11432_/Q _05914_/A2 _06806_/B1 _10505_/Q vssd1 vssd1 vccd1 vccd1 _05914_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_95_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ _09692_/B _09682_/B vssd1 vssd1 vccd1 vccd1 _09682_/Y sky130_fd_sc_hd__nand2_2
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06894_ _10216_/Q _09959_/A vssd1 vssd1 vccd1 vccd1 _08243_/D sky130_fd_sc_hd__nand2_2
XFILLER_82_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08633_ _11171_/Q _08633_/B vssd1 vssd1 vccd1 vccd1 _08633_/X sky130_fd_sc_hd__or2_1
X_05845_ _10266_/Q _06998_/A _06373_/B1 _10311_/Q vssd1 vssd1 vccd1 vccd1 _05845_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _08745_/A _08577_/S vssd1 vssd1 vccd1 vccd1 _08901_/S sky130_fd_sc_hd__or2_4
XFILLER_23_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05776_ _10507_/Q _06998_/A _07111_/A _10310_/Q vssd1 vssd1 vccd1 vccd1 _05776_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07515_ input92/X _10542_/Q _07533_/S vssd1 vssd1 vccd1 vccd1 _07516_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08495_ _08970_/A1 _11098_/Q _08501_/S vssd1 vssd1 vccd1 vccd1 _08496_/B sky130_fd_sc_hd__mux2_1
XFILLER_74_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07446_ _07785_/A0 _07513_/S _07442_/Y _10498_/Q _09193_/A vssd1 vssd1 vccd1 vccd1
+ _10498_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07377_ _10463_/Q _07010_/A _07393_/S vssd1 vssd1 vccd1 vccd1 _07378_/B sky130_fd_sc_hd__mux2_1
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09116_ _10165_/A1 _09110_/X _09115_/X _09279_/C1 vssd1 vssd1 vccd1 vccd1 _11404_/D
+ sky130_fd_sc_hd__o211a_1
X_06328_ _10881_/Q _06468_/B _06152_/B _10929_/Q _07083_/B vssd1 vssd1 vccd1 vccd1
+ _06328_/X sky130_fd_sc_hd__o221a_1
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09047_ _11373_/Q _09055_/B vssd1 vssd1 vccd1 vccd1 _09047_/X sky130_fd_sc_hd__or2_1
X_06259_ _11262_/Q _06635_/B1 _06126_/B _11214_/Q _06258_/X vssd1 vssd1 vccd1 vccd1
+ _06259_/X sky130_fd_sc_hd__o221a_1
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout930 input99/X vssd1 vssd1 vccd1 vccd1 _07002_/A sky130_fd_sc_hd__buf_6
Xfanout941 input96/X vssd1 vssd1 vccd1 vccd1 _09237_/A0 sky130_fd_sc_hd__clkbuf_16
X_09949_ _10372_/Q _09570_/A _09570_/B _10692_/Q vssd1 vssd1 vccd1 vccd1 _09949_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout952 fanout958/X vssd1 vssd1 vccd1 vccd1 _08838_/A0 sky130_fd_sc_hd__clkbuf_8
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout963 _07104_/A vssd1 vssd1 vccd1 vccd1 _10132_/A0 sky130_fd_sc_hd__buf_6
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout974 _08929_/A1 vssd1 vssd1 vccd1 vccd1 _08876_/A0 sky130_fd_sc_hd__buf_6
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout985 input84/X vssd1 vssd1 vccd1 vccd1 _11871_/A sky130_fd_sc_hd__buf_8
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout996 _06849_/C1 vssd1 vssd1 vccd1 vccd1 _06997_/A sky130_fd_sc_hd__buf_6
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1087 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1087/HI io_oeb[17] sky130_fd_sc_hd__conb_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1098 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1098/HI io_oeb[28] sky130_fd_sc_hd__conb_1
X_11773_ _11781_/CLK _11773_/D vssd1 vssd1 vccd1 vccd1 _11773_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _10798_/CLK _10724_/D vssd1 vssd1 vccd1 vccd1 _10724_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10655_ _10805_/CLK _10655_/D vssd1 vssd1 vccd1 vccd1 _10655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10586_ _11628_/CLK _10586_/D vssd1 vssd1 vccd1 vccd1 _10586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ _11325_/CLK _11207_/D vssd1 vssd1 vccd1 vccd1 _11207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11138_ _11224_/CLK _11138_/D vssd1 vssd1 vccd1 vccd1 _11138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11069_ _11766_/CLK _11069_/D vssd1 vssd1 vccd1 vccd1 _11069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05630_ _11785_/Q _05630_/A2 _05630_/B1 _11783_/Q _05628_/X vssd1 vssd1 vccd1 vccd1
+ _05633_/A sky130_fd_sc_hd__a221o_4
XFILLER_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05561_ _05561_/A _05561_/B vssd1 vssd1 vccd1 vccd1 _05561_/Y sky130_fd_sc_hd__nor2_8
XFILLER_60_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07300_ _07300_/A _08665_/C _10087_/C vssd1 vssd1 vccd1 vccd1 _08760_/S sky130_fd_sc_hd__or3_4
X_05492_ _10237_/Q input48/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05492_/X sky130_fd_sc_hd__mux2_2
X_08280_ _10972_/Q _08284_/B vssd1 vssd1 vccd1 vccd1 _08280_/X sky130_fd_sc_hd__or2_1
XFILLER_32_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07231_ _07095_/X _10383_/Q _07233_/S vssd1 vssd1 vccd1 vccd1 _10383_/D sky130_fd_sc_hd__mux2_1
X_07162_ _10017_/A0 _10342_/Q _09243_/C vssd1 vssd1 vccd1 vccd1 _07163_/B sky130_fd_sc_hd__mux2_1
XFILLER_34_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06113_ _11464_/Q _07152_/A _06112_/X _06808_/C1 vssd1 vssd1 vccd1 vccd1 _06113_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07093_ _07318_/A _07229_/B vssd1 vssd1 vccd1 vccd1 _07093_/X sky130_fd_sc_hd__or2_4
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06044_ _10750_/Q _07853_/A _07455_/A _10657_/Q vssd1 vssd1 vccd1 vccd1 _06044_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout215 _07820_/Y vssd1 vssd1 vccd1 vccd1 _07959_/S sky130_fd_sc_hd__buf_6
XFILLER_99_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout226 _07205_/Y vssd1 vssd1 vccd1 vccd1 _07772_/S sky130_fd_sc_hd__buf_4
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09803_ _10288_/Q _09573_/B _09573_/C _10296_/Q vssd1 vssd1 vccd1 vccd1 _09803_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout237 _10025_/S vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_101_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout248 _08874_/S vssd1 vssd1 vccd1 vccd1 _08890_/S sky130_fd_sc_hd__buf_6
Xfanout259 _08567_/S vssd1 vssd1 vccd1 vccd1 _08577_/S sky130_fd_sc_hd__buf_6
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07995_ _10822_/Q _08091_/C vssd1 vssd1 vccd1 vccd1 _07995_/X sky130_fd_sc_hd__or2_1
XFILLER_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09734_ _10341_/Q _09886_/A2 _09881_/B1 _11465_/Q _09733_/X vssd1 vssd1 vccd1 vccd1
+ _09739_/B sky130_fd_sc_hd__a221o_1
XFILLER_101_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06946_ _09431_/B _06945_/X _06942_/A vssd1 vssd1 vccd1 vccd1 _06969_/S sky130_fd_sc_hd__a21o_4
XFILLER_55_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10939_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09665_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _11631_/D sky130_fd_sc_hd__nand2_1
X_06877_ _11477_/Q _07153_/A _06877_/B1 _11401_/Q _06876_/X vssd1 vssd1 vccd1 vccd1
+ _06877_/X sky130_fd_sc_hd__o221a_1
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08616_ _08876_/A0 _08623_/S _08615_/X _08947_/C1 vssd1 vssd1 vccd1 vccd1 _11162_/D
+ sky130_fd_sc_hd__o211a_1
X_05828_ _11489_/Q _08907_/A _08855_/A _11413_/Q _06670_/D1 vssd1 vssd1 vccd1 vccd1
+ _05828_/X sky130_fd_sc_hd__o221a_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _09594_/X _09596_/B vssd1 vssd1 vccd1 vccd1 _09817_/B sky130_fd_sc_hd__nand2b_1
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _11123_/Q _07353_/B _07355_/S _07324_/B vssd1 vssd1 vccd1 vccd1 _11123_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05759_ _11369_/Q _06221_/A2 _09110_/A _11402_/Q _05758_/X vssd1 vssd1 vccd1 vccd1
+ _05759_/X sky130_fd_sc_hd__o221a_2
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08478_ _08579_/A0 _08501_/S _08477_/X _09036_/C1 vssd1 vssd1 vccd1 vccd1 _11089_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07429_ _07034_/A _10491_/Q _07429_/S vssd1 vssd1 vccd1 vccd1 _07430_/B sky130_fd_sc_hd__mux2_1
XFILLER_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10440_ _11177_/CLK _10440_/D vssd1 vssd1 vccd1 vccd1 _10440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10371_ _11713_/CLK _10371_/D vssd1 vssd1 vccd1 vccd1 _10371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout760 _06674_/A2 vssd1 vssd1 vccd1 vccd1 _06806_/B1 sky130_fd_sc_hd__buf_2
XFILLER_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout771 fanout782/X vssd1 vssd1 vccd1 vccd1 _10119_/A sky130_fd_sc_hd__buf_6
Xfanout782 fanout793/X vssd1 vssd1 vccd1 vccd1 fanout782/X sky130_fd_sc_hd__buf_6
XFILLER_120_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout793 _05747_/Y vssd1 vssd1 vccd1 vccd1 fanout793/X sky130_fd_sc_hd__buf_12
XFILLER_150_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _10134_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _10023_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 _05434_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _07052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_164 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_175 fanout738/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 _08818_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _10021_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11756_ _11756_/CLK _11756_/D vssd1 vssd1 vccd1 vccd1 _11756_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10707_ _11573_/CLK _10707_/D vssd1 vssd1 vccd1 vccd1 _10707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11687_ _11735_/CLK _11687_/D vssd1 vssd1 vccd1 vccd1 _11687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10638_ _11270_/CLK _10638_/D vssd1 vssd1 vccd1 vccd1 _10638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10569_ _10769_/CLK _10569_/D vssd1 vssd1 vccd1 vccd1 _10569_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06800_ _10629_/Q _06871_/A2 _07539_/A _10355_/Q vssd1 vssd1 vccd1 vccd1 _06800_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07780_ _07796_/A _07780_/B vssd1 vssd1 vccd1 vccd1 _10697_/D sky130_fd_sc_hd__or2_1
XFILLER_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 io_in[8] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
X_06731_ _10693_/Q _07202_/A _06731_/B1 _10516_/Q _06725_/X vssd1 vssd1 vccd1 vccd1
+ _06731_/X sky130_fd_sc_hd__o221a_1
XFILLER_83_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09450_ _09441_/B input11/X _09441_/Y input28/X _09449_/X vssd1 vssd1 vccd1 vccd1
+ _09450_/X sky130_fd_sc_hd__a221o_1
XFILLER_92_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06662_ _07081_/A _06633_/X _06644_/X _06661_/X vssd1 vssd1 vccd1 vccd1 _06662_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_65_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08401_ _08847_/A _08401_/B vssd1 vssd1 vccd1 vccd1 _11041_/D sky130_fd_sc_hd__or2_1
X_05613_ _05075_/Y _11398_/Q _11394_/Q _05077_/Y _05610_/X vssd1 vssd1 vccd1 vccd1
+ _05613_/X sky130_fd_sc_hd__a221o_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09381_ _09999_/A0 _11548_/Q _09390_/S vssd1 vssd1 vccd1 vccd1 _11548_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06593_ _10741_/Q _06634_/B1 _07111_/A _11780_/Q _06592_/X vssd1 vssd1 vccd1 vccd1
+ _06593_/X sky130_fd_sc_hd__o221a_1
XFILLER_80_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08332_ _11007_/Q _08322_/Y _08325_/Y _07316_/X vssd1 vssd1 vccd1 vccd1 _11007_/D
+ sky130_fd_sc_hd__a22o_1
X_05544_ _05616_/A1 _11495_/Q _11492_/Q _05077_/A vssd1 vssd1 vccd1 vccd1 _05544_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08263_ _08793_/A _08263_/B vssd1 vssd1 vccd1 vccd1 _10963_/D sky130_fd_sc_hd__or2_1
XFILLER_20_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05475_ _11604_/Q _11603_/Q _09477_/A _05475_/D vssd1 vssd1 vccd1 vccd1 _05475_/X
+ sky130_fd_sc_hd__and4b_4
X_07214_ _07031_/A _07205_/B _07772_/S _10371_/Q vssd1 vssd1 vccd1 vccd1 _10371_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08194_ _10932_/Q _08197_/S _07644_/Y _08817_/B2 vssd1 vssd1 vccd1 vccd1 _10932_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_69_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07145_ _10334_/Q _07145_/B vssd1 vssd1 vccd1 vccd1 _07145_/X sky130_fd_sc_hd__or2_1
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07076_ _07076_/A _07205_/A vssd1 vssd1 vccd1 vccd1 _07187_/B sky130_fd_sc_hd__and2_4
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06027_ _11426_/Q _09154_/A _06026_/X _06670_/D1 vssd1 vssd1 vccd1 vccd1 _06027_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07978_ _08733_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _10812_/D sky130_fd_sc_hd__or2_1
X_09717_ _10398_/Q _09873_/A2 _09875_/A2 _11432_/Q vssd1 vssd1 vccd1 vccd1 _09717_/X
+ sky130_fd_sc_hd__a22o_1
X_06929_ _10185_/A0 _10207_/Q _06934_/S vssd1 vssd1 vccd1 vccd1 _10207_/D sky130_fd_sc_hd__mux2_1
X_09648_ _10323_/Q _09948_/B1 _09947_/B1 _10328_/Q vssd1 vssd1 vccd1 vccd1 _09648_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _10270_/Q _09571_/B _09573_/D _10269_/Q vssd1 vssd1 vccd1 vccd1 _09579_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11610_ _11663_/CLK _11610_/D vssd1 vssd1 vccd1 vccd1 _11610_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11541_ _11801_/CLK _11541_/D vssd1 vssd1 vccd1 vccd1 _11541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11472_ _11472_/CLK _11472_/D vssd1 vssd1 vccd1 vccd1 _11472_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_137_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10423_ _11233_/CLK _10423_/D vssd1 vssd1 vccd1 vccd1 _10423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10354_ _10798_/CLK _10354_/D vssd1 vssd1 vccd1 vccd1 _10354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10285_ _10812_/CLK _10285_/D vssd1 vssd1 vccd1 vccd1 _10285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout590 _06743_/A vssd1 vssd1 vccd1 vccd1 _06855_/B sky130_fd_sc_hd__buf_12
XFILLER_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _11808_/CLK _11808_/D vssd1 vssd1 vccd1 vccd1 _11808_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11739_ _11762_/CLK _11739_/D vssd1 vssd1 vccd1 vccd1 _11739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05260_ _10442_/Q _10441_/Q _05392_/S vssd1 vssd1 vccd1 vccd1 _05264_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05191_ _05413_/S _11065_/Q vssd1 vssd1 vccd1 vccd1 _05191_/X sky130_fd_sc_hd__and2_1
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08950_ _11602_/Q _08950_/B vssd1 vssd1 vccd1 vccd1 _09554_/A sky130_fd_sc_hd__nand2_4
XFILLER_142_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07901_ _10769_/Q _07901_/B vssd1 vssd1 vccd1 vccd1 _07901_/X sky130_fd_sc_hd__or2_1
X_08881_ _08941_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _11297_/D sky130_fd_sc_hd__or2_1
XFILLER_97_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07832_ _10134_/A0 _07820_/B _07821_/A _10727_/Q vssd1 vssd1 vccd1 vccd1 _10727_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07763_ _10683_/Q _07008_/X _07772_/S vssd1 vssd1 vccd1 vccd1 _10683_/D sky130_fd_sc_hd__mux2_1
X_09502_ _09502_/A _09502_/B _09500_/C vssd1 vssd1 vccd1 vccd1 _09502_/X sky130_fd_sc_hd__or3b_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06714_ _10275_/Q _06858_/B1 _06711_/X _06713_/X _06997_/A vssd1 vssd1 vccd1 vccd1
+ _06714_/X sky130_fd_sc_hd__o2111a_1
XFILLER_77_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07694_ _08323_/A _08589_/S vssd1 vssd1 vccd1 vccd1 _07694_/Y sky130_fd_sc_hd__nand2_2
XFILLER_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09433_ _11629_/Q _09692_/B vssd1 vssd1 vccd1 vccd1 _09434_/B sky130_fd_sc_hd__nor2_1
X_06645_ _10406_/Q _06645_/A2 _08971_/A _10569_/Q vssd1 vssd1 vccd1 vccd1 _06645_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09364_ _09364_/A1 _09376_/B _10156_/B1 vssd1 vssd1 vccd1 vccd1 _09364_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06576_ _06576_/A _06576_/B _06576_/C vssd1 vssd1 vccd1 vccd1 _06576_/X sky130_fd_sc_hd__or3_1
X_08315_ _10112_/A0 _10994_/Q _08321_/S vssd1 vssd1 vccd1 vccd1 _10994_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05527_ _11628_/Q _11506_/Q _11500_/Q _11625_/Q vssd1 vssd1 vccd1 vccd1 _05527_/X
+ sky130_fd_sc_hd__a22o_1
X_09295_ _11498_/Q _09293_/X _09294_/X vssd1 vssd1 vccd1 vccd1 _11498_/D sky130_fd_sc_hd__a21o_1
XANTENNA_20 _06558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 _07022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_42 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _10955_/Q _08284_/B vssd1 vssd1 vccd1 vccd1 _08246_/X sky130_fd_sc_hd__or2_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_64 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05458_ _10754_/Q _09947_/A2 _09873_/A2 _10750_/Q vssd1 vssd1 vccd1 vccd1 _05458_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_75 _11614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_86 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_97 _09572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ _07059_/A _10919_/Q _08181_/S vssd1 vssd1 vccd1 vccd1 _10919_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05389_ _05389_/A _05389_/B _05389_/C _05389_/D vssd1 vssd1 vccd1 vccd1 _05390_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_107_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07128_ _10324_/Q _07145_/B vssd1 vssd1 vccd1 vccd1 _07128_/X sky130_fd_sc_hd__or2_1
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07059_ _07059_/A _10028_/A vssd1 vssd1 vccd1 vccd1 _07316_/B sky130_fd_sc_hd__and2_4
Xoutput160 _11580_/Q vssd1 vssd1 vccd1 vccd1 rom_addr[2] sky130_fd_sc_hd__buf_4
XFILLER_0_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput171 _11869_/X vssd1 vssd1 vccd1 vccd1 wb_rom_adrb[3] sky130_fd_sc_hd__buf_4
XFILLER_88_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput182 _05488_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_4
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10070_ _10117_/A0 _11731_/Q _10071_/S vssd1 vssd1 vccd1 vccd1 _11731_/D sky130_fd_sc_hd__mux2_1
Xoutput193 _05498_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_4
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10972_ _11812_/CLK _10972_/D vssd1 vssd1 vccd1 vccd1 _10972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11524_ _11527_/CLK _11524_/D vssd1 vssd1 vccd1 vccd1 _11524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11455_ _11644_/CLK _11455_/D vssd1 vssd1 vccd1 vccd1 _11455_/Q sky130_fd_sc_hd__dfxtp_1
X_10406_ _10769_/CLK _10406_/D vssd1 vssd1 vccd1 vccd1 _10406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11386_ _11683_/CLK _11386_/D vssd1 vssd1 vccd1 vccd1 _11386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10337_ _11471_/CLK _10337_/D vssd1 vssd1 vccd1 vccd1 _10337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _11713_/CLK _10268_/D vssd1 vssd1 vccd1 vccd1 _10268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10199_ _11803_/CLK _10199_/D vssd1 vssd1 vccd1 vccd1 _10199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06430_ _10848_/Q _06430_/A2 _06426_/X _06429_/X vssd1 vssd1 vccd1 vccd1 _06431_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06361_ _11791_/Q _09132_/A _09293_/A _11507_/Q _06360_/X vssd1 vssd1 vccd1 vccd1
+ _06361_/X sky130_fd_sc_hd__o221a_1
XFILLER_148_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08100_ _10874_/Q _08437_/A _08354_/S _08303_/A vssd1 vssd1 vccd1 vccd1 _08100_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_72_1288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05312_ _05312_/A _05312_/B _05312_/C _05312_/D vssd1 vssd1 vccd1 vccd1 _05313_/B
+ sky130_fd_sc_hd__or4_4
X_09080_ _11388_/Q _09060_/X _09079_/X vssd1 vssd1 vccd1 vccd1 _11388_/D sky130_fd_sc_hd__a21o_1
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06292_ _11387_/Q _09060_/A _08668_/A _11430_/Q _06291_/X vssd1 vssd1 vccd1 vccd1
+ _06292_/X sky130_fd_sc_hd__o221a_1
XFILLER_30_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08031_ _08876_/A0 _10840_/Q _08035_/S vssd1 vssd1 vccd1 vccd1 _08032_/B sky130_fd_sc_hd__mux2_1
Xinput40 rom_value[8] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_2
X_05243_ _09539_/B _10861_/Q _10790_/Q _05414_/S vssd1 vssd1 vccd1 vccd1 _05247_/A
+ sky130_fd_sc_hd__a22o_1
Xinput51 wb_rom_val[18] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_4
Xinput62 wb_rom_val[28] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_4
Xinput73 wb_rom_val[9] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__buf_2
XFILLER_115_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput84 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_4
Xinput95 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__buf_4
X_05174_ _11226_/Q _11225_/Q _05377_/S vssd1 vssd1 vccd1 vccd1 _05176_/C sky130_fd_sc_hd__mux2_1
XFILLER_143_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09982_ _10165_/A1 _09994_/B _10178_/B1 vssd1 vssd1 vccd1 vccd1 _09982_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08933_ _08933_/A1 _08940_/S _08932_/X _08943_/C1 vssd1 vssd1 vccd1 vccd1 _11325_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08864_ _11289_/Q _08894_/B vssd1 vssd1 vccd1 vccd1 _08864_/X sky130_fd_sc_hd__or2_1
XFILLER_97_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07815_ input103/X _10715_/Q _07817_/S vssd1 vssd1 vccd1 vccd1 _07816_/B sky130_fd_sc_hd__mux2_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08795_ _08937_/A1 _08792_/S _08794_/X _08937_/C1 vssd1 vssd1 vccd1 vccd1 _11253_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07746_ _10674_/Q _07760_/B vssd1 vssd1 vccd1 vccd1 _07746_/X sky130_fd_sc_hd__or2_1
XFILLER_84_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07677_ _10633_/Q _07673_/Y _07676_/X _08440_/B2 vssd1 vssd1 vccd1 vccd1 _10633_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09416_ _09416_/A _09416_/B vssd1 vssd1 vccd1 vccd1 _09426_/S sky130_fd_sc_hd__nand2_4
XFILLER_52_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06628_ _10833_/Q _07994_/A _06628_/B1 _11278_/Q vssd1 vssd1 vccd1 vccd1 _06628_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09347_ _09347_/A _10108_/B _10119_/C vssd1 vssd1 vccd1 vccd1 _09357_/S sky130_fd_sc_hd__or3_4
X_06559_ _06546_/X _06547_/X _06558_/X _06619_/A1 vssd1 vssd1 vccd1 vccd1 _06576_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09278_ _11491_/Q _09288_/B vssd1 vssd1 vccd1 vccd1 _09278_/X sky130_fd_sc_hd__or2_1
XFILLER_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08229_ _08560_/A _08471_/B _10136_/C vssd1 vssd1 vccd1 vccd1 _08324_/B sky130_fd_sc_hd__and3_4
XFILLER_153_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11240_ _11393_/CLK _11240_/D vssd1 vssd1 vccd1 vccd1 _11240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11171_ _11812_/CLK _11171_/D vssd1 vssd1 vccd1 vccd1 _11171_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_122_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10122_ _07007_/A _11768_/Q _10134_/S vssd1 vssd1 vccd1 vccd1 _11768_/D sky130_fd_sc_hd__mux2_1
X_10053_ _11718_/Q _07141_/A _10057_/S vssd1 vssd1 vccd1 vccd1 _10054_/B sky130_fd_sc_hd__mux2_1
XFILLER_76_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10955_ _11291_/CLK _10955_/D vssd1 vssd1 vccd1 vccd1 _10955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10886_ _10929_/CLK _10886_/D vssd1 vssd1 vccd1 vccd1 _10886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11507_ _11800_/CLK _11507_/D vssd1 vssd1 vccd1 vccd1 _11507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11438_ _11473_/CLK _11438_/D vssd1 vssd1 vccd1 vccd1 _11438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11369_ _11495_/CLK _11369_/D vssd1 vssd1 vccd1 vccd1 _11369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05930_ _10603_/Q _06635_/B1 _06636_/A2 _11071_/Q vssd1 vssd1 vccd1 vccd1 _05930_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05861_ _11182_/Q _08650_/A _10119_/A _10452_/Q vssd1 vssd1 vccd1 vccd1 _05864_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07600_ _09229_/A _08850_/S vssd1 vssd1 vccd1 vccd1 _07600_/Y sky130_fd_sc_hd__nand2_2
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08580_ _08833_/A _08580_/B vssd1 vssd1 vccd1 vccd1 _11145_/D sky130_fd_sc_hd__or2_1
XFILLER_130_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05792_ _11103_/Q _06716_/A2 _05789_/Y _05791_/X vssd1 vssd1 vccd1 vccd1 _05792_/X
+ sky130_fd_sc_hd__o211a_1
X_07531_ _07141_/A _10550_/Q _07533_/S vssd1 vssd1 vccd1 vccd1 _07532_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07462_ _10026_/A _07462_/B vssd1 vssd1 vccd1 vccd1 _10508_/D sky130_fd_sc_hd__or2_1
XFILLER_90_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09201_ _09201_/A1 _09200_/X _07441_/A vssd1 vssd1 vccd1 vccd1 _11447_/D sky130_fd_sc_hd__a21o_1
X_06413_ _11065_/Q _06413_/A2 _06411_/X _06412_/X vssd1 vssd1 vccd1 vccd1 _06413_/X
+ sky130_fd_sc_hd__o211a_1
X_07393_ _10473_/Q _10135_/A0 _07393_/S vssd1 vssd1 vccd1 vccd1 _07394_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_56_wb_clk_i clkbuf_leaf_88_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11628_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09132_ _09132_/A _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09132_/X sky130_fd_sc_hd__or3_4
X_06344_ _11695_/Q _09998_/A _06924_/A _11742_/Q _06344_/C1 vssd1 vssd1 vccd1 vccd1
+ _06344_/X sky130_fd_sc_hd__o221a_1
XFILLER_108_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09063_ _11380_/Q _09077_/B vssd1 vssd1 vccd1 vccd1 _09063_/X sky130_fd_sc_hd__or2_1
XFILLER_11_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06275_ _05816_/A _06212_/Y _05820_/B vssd1 vssd1 vccd1 vccd1 _06275_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08014_ _07107_/A _08011_/S _08013_/X _08841_/C1 vssd1 vssd1 vccd1 vccd1 _10831_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05226_ _10951_/Q _11003_/Q _05416_/S vssd1 vssd1 vccd1 vccd1 _05237_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05157_ _05157_/A _05157_/B vssd1 vssd1 vccd1 vccd1 _05157_/Y sky130_fd_sc_hd__nor2_8
XFILLER_131_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09965_ _09965_/A _10108_/B _10119_/C vssd1 vssd1 vccd1 vccd1 _09975_/S sky130_fd_sc_hd__or3_4
X_05088_ _05427_/S vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__inv_4
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08916_ _11317_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08916_/X sky130_fd_sc_hd__or2_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _11699_/Q _09568_/B _09947_/B1 _11714_/Q _09895_/X vssd1 vssd1 vccd1 vccd1
+ _09899_/C sky130_fd_sc_hd__a221o_1
XFILLER_57_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _08847_/A _08847_/B vssd1 vssd1 vccd1 vccd1 _11281_/D sky130_fd_sc_hd__or2_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08778_ _11245_/Q _08804_/B vssd1 vssd1 vccd1 vccd1 _08778_/X sky130_fd_sc_hd__or2_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _08846_/A0 _07761_/A2 _07728_/X _07902_/C1 vssd1 vssd1 vccd1 vccd1 _10665_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_26_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10740_ _11780_/CLK _10740_/D vssd1 vssd1 vccd1 vccd1 _10740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _10785_/CLK _10671_/D vssd1 vssd1 vccd1 vccd1 _10671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11223_ _11307_/CLK _11223_/D vssd1 vssd1 vccd1 vccd1 _11223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ _11527_/CLK _11154_/D vssd1 vssd1 vccd1 vccd1 _11154_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10105_ _10105_/A1 _10087_/X _10104_/X _10155_/C1 vssd1 vssd1 vccd1 vccd1 _11754_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11085_ _11651_/CLK _11085_/D vssd1 vssd1 vccd1 vccd1 _11085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10036_ _11708_/Q _08661_/A _10051_/S vssd1 vssd1 vccd1 vccd1 _10037_/B sky130_fd_sc_hd__mux2_1
XFILLER_76_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10938_ _11756_/CLK _10938_/D vssd1 vssd1 vccd1 vccd1 _10938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10869_ _11270_/CLK _10869_/D vssd1 vssd1 vccd1 vccd1 _10869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06060_ _10459_/Q _06308_/A2 _06373_/B1 _10812_/Q vssd1 vssd1 vccd1 vccd1 _06060_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout408 _05379_/Y vssd1 vssd1 vccd1 vccd1 _09948_/B1 sky130_fd_sc_hd__buf_8
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout419 _05324_/Y vssd1 vssd1 vccd1 vccd1 _09878_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_103_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11470_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09750_ _10549_/Q _09882_/B1 _09567_/D _10544_/Q vssd1 vssd1 vccd1 vccd1 _09750_/X
+ sky130_fd_sc_hd__a22o_1
X_06962_ _06967_/A _06961_/X _06969_/S vssd1 vssd1 vccd1 vccd1 _06962_/X sky130_fd_sc_hd__mux2_4
XFILLER_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05913_ _10748_/Q _06861_/B _06806_/A2 _10556_/Q vssd1 vssd1 vccd1 vccd1 _05913_/X
+ sky130_fd_sc_hd__o22a_1
X_08701_ _11205_/Q _08705_/B vssd1 vssd1 vccd1 vccd1 _08701_/X sky130_fd_sc_hd__or2_1
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09681_ _09681_/A _09681_/B _09681_/C _09681_/D vssd1 vssd1 vccd1 vccd1 _09682_/B
+ sky130_fd_sc_hd__or4_4
X_06893_ _10216_/Q _09959_/A vssd1 vssd1 vccd1 vccd1 _07151_/D sky130_fd_sc_hd__and2_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08632_ _08893_/A1 _08623_/S _08631_/X _09078_/C1 vssd1 vssd1 vccd1 vccd1 _11170_/D
+ sky130_fd_sc_hd__o211a_1
X_05844_ _10380_/Q _06371_/A2 _06105_/B1 _10795_/Q vssd1 vssd1 vccd1 vccd1 _05844_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08563_ _08745_/A _08577_/S vssd1 vssd1 vccd1 vccd1 _08563_/Y sky130_fd_sc_hd__nor2_2
X_05775_ _10379_/Q _07222_/A _07819_/A _10717_/Q vssd1 vssd1 vccd1 vccd1 _05775_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07514_ _07916_/A _07514_/B vssd1 vssd1 vccd1 vccd1 _10541_/D sky130_fd_sc_hd__or2_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08494_ _08969_/A1 _08501_/S _08493_/X _08662_/C1 vssd1 vssd1 vccd1 vccd1 _11097_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07445_ _10015_/A0 _07513_/S _07442_/Y _10497_/Q _09193_/A vssd1 vssd1 vccd1 vccd1
+ _10497_/D sky130_fd_sc_hd__o221a_1
XFILLER_126_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07376_ _10462_/Q _07380_/S _07655_/S _07090_/A vssd1 vssd1 vccd1 vccd1 _10462_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09115_ _11404_/Q _09127_/B vssd1 vssd1 vccd1 vccd1 _09115_/X sky130_fd_sc_hd__or2_1
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06327_ _10853_/Q _06631_/A2 _06323_/X _06326_/X vssd1 vssd1 vccd1 vccd1 _06327_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09046_ _09090_/A1 _09038_/X _09045_/X _09289_/C1 vssd1 vssd1 vccd1 vccd1 _11372_/D
+ sky130_fd_sc_hd__o211a_1
X_06258_ _10442_/Q _06513_/A2 _08647_/B _11178_/Q vssd1 vssd1 vccd1 vccd1 _06258_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05209_ _09538_/A _10904_/Q _10427_/Q _09539_/B vssd1 vssd1 vccd1 vccd1 _05213_/A
+ sky130_fd_sc_hd__a22o_1
X_06189_ _06189_/A1 _06183_/X _06188_/X _08243_/A _06178_/X vssd1 vssd1 vccd1 vccd1
+ _06189_/X sky130_fd_sc_hd__o311a_2
XFILLER_117_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout920 _06297_/C1 vssd1 vssd1 vccd1 vccd1 _06651_/C1 sky130_fd_sc_hd__buf_6
XFILLER_89_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout931 _09114_/A1 vssd1 vssd1 vccd1 vccd1 _09275_/A1 sky130_fd_sc_hd__buf_6
Xfanout942 _09216_/A0 vssd1 vssd1 vccd1 vccd1 _07025_/A sky130_fd_sc_hd__buf_6
X_09948_ _10690_/Q _09565_/B _09948_/B1 _10368_/Q _09947_/X vssd1 vssd1 vccd1 vccd1
+ _09957_/C sky130_fd_sc_hd__a221o_1
Xfanout953 fanout958/X vssd1 vssd1 vccd1 vccd1 _10134_/A0 sky130_fd_sc_hd__buf_8
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout964 _07104_/A vssd1 vssd1 vccd1 vccd1 _08834_/A0 sky130_fd_sc_hd__buf_4
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout975 input89/X vssd1 vssd1 vccd1 vccd1 _08929_/A1 sky130_fd_sc_hd__clkbuf_16
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout986 _07689_/A vssd1 vssd1 vccd1 vccd1 _06633_/A sky130_fd_sc_hd__buf_4
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _10580_/Q _09879_/A2 _09879_/B1 _10574_/Q _09878_/X vssd1 vssd1 vccd1 vccd1
+ _09880_/D sky130_fd_sc_hd__a221o_4
Xfanout997 _06670_/D1 vssd1 vssd1 vccd1 vccd1 _06849_/C1 sky130_fd_sc_hd__buf_6
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1088 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1088/HI io_oeb[18] sky130_fd_sc_hd__conb_1
XFILLER_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11772_ _11776_/CLK _11772_/D vssd1 vssd1 vccd1 vccd1 _11772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1099 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1099/HI io_oeb[29] sky130_fd_sc_hd__conb_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10723_ _10727_/CLK _10723_/D vssd1 vssd1 vccd1 vccd1 _10723_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10654_ _10765_/CLK _10654_/D vssd1 vssd1 vccd1 vccd1 _10654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10585_ _11280_/CLK _10585_/D vssd1 vssd1 vccd1 vccd1 _10585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11770_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11206_ _11812_/CLK _11206_/D vssd1 vssd1 vccd1 vccd1 _11206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11137_ _11224_/CLK _11137_/D vssd1 vssd1 vccd1 vccd1 _11137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11068_ _11186_/CLK _11068_/D vssd1 vssd1 vccd1 vccd1 _11068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10019_ _10019_/A0 _11700_/Q _10028_/B vssd1 vssd1 vccd1 vccd1 _10020_/B sky130_fd_sc_hd__mux2_1
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05560_ _05076_/A _11345_/Q _11340_/Q _05620_/B2 _05559_/X vssd1 vssd1 vccd1 vccd1
+ _05561_/B sky130_fd_sc_hd__a221o_4
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05491_ _10236_/Q input47/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05491_/X sky130_fd_sc_hd__mux2_2
XFILLER_60_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07230_ _07229_/X _10382_/Q _07233_/S vssd1 vssd1 vccd1 vccd1 _10382_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07161_ _07920_/A _07161_/B vssd1 vssd1 vccd1 vccd1 _10341_/D sky130_fd_sc_hd__or2_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06112_ _10702_/Q _07778_/A _07853_/A _10804_/Q _06111_/X vssd1 vssd1 vccd1 vccd1
+ _06112_/X sky130_fd_sc_hd__o221a_2
X_07092_ _07092_/A _10028_/A vssd1 vssd1 vccd1 vccd1 _07229_/B sky130_fd_sc_hd__and2_4
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06043_ _10478_/Q _06803_/A2 _06857_/B1 _11699_/Q _06997_/A vssd1 vssd1 vccd1 vccd1
+ _06043_/X sky130_fd_sc_hd__o221a_1
XFILLER_126_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout216 _07624_/Y vssd1 vssd1 vccd1 vccd1 _07628_/S sky130_fd_sc_hd__buf_4
Xfanout227 _07204_/Y vssd1 vssd1 vccd1 vccd1 _07771_/B1 sky130_fd_sc_hd__buf_8
X_09802_ _10285_/Q _09571_/B _09572_/D _10286_/Q vssd1 vssd1 vccd1 vccd1 _09802_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout238 _10009_/Y vssd1 vssd1 vccd1 vccd1 _10051_/S sky130_fd_sc_hd__buf_6
X_07994_ _07994_/A _08665_/C _09038_/C vssd1 vssd1 vccd1 vccd1 _07994_/X sky130_fd_sc_hd__or3_4
Xfanout249 _08874_/S vssd1 vssd1 vccd1 vccd1 _08884_/S sky130_fd_sc_hd__buf_2
XFILLER_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09733_ _11475_/Q _09871_/A2 _09877_/B1 _11466_/Q _09732_/X vssd1 vssd1 vccd1 vccd1
+ _09733_/X sky130_fd_sc_hd__a221o_1
X_06945_ _11599_/Q _06945_/B _09538_/A vssd1 vssd1 vccd1 vccd1 _06945_/X sky130_fd_sc_hd__or3_1
XFILLER_132_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06876_ _11440_/Q _07254_/A _07440_/A _10553_/Q vssd1 vssd1 vccd1 vccd1 _06876_/X
+ sky130_fd_sc_hd__o22a_1
X_09664_ _11631_/Q _09959_/B _09959_/A vssd1 vssd1 vccd1 vccd1 _09665_/B sky130_fd_sc_hd__a21oi_1
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05827_ _11423_/Q _08668_/A _09038_/A _11370_/Q vssd1 vssd1 vccd1 vccd1 _05827_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08615_ _11162_/Q _08633_/B vssd1 vssd1 vccd1 vccd1 _08615_/X sky130_fd_sc_hd__or2_1
X_09595_ _09594_/B _09594_/C _09594_/D _11658_/Q vssd1 vssd1 vccd1 vccd1 _09596_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_83_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11410_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05758_ _11488_/Q _09271_/A _06717_/B1 _11339_/Q vssd1 vssd1 vccd1 vccd1 _05758_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08546_ _08947_/A1 _08529_/S _08545_/X _08921_/C1 vssd1 vssd1 vccd1 vccd1 _11122_/D
+ sky130_fd_sc_hd__o211a_1
X_08477_ _11089_/Q _08503_/B vssd1 vssd1 vccd1 vccd1 _08477_/X sky130_fd_sc_hd__or2_1
X_05689_ _11171_/Q _05518_/Y _05621_/Y _11164_/Q vssd1 vssd1 vccd1 vccd1 _05689_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07428_ _10043_/A _07428_/B vssd1 vssd1 vccd1 vccd1 _10490_/D sky130_fd_sc_hd__or2_1
XFILLER_52_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07359_ _08196_/A _07991_/S vssd1 vssd1 vccd1 vccd1 _07363_/S sky130_fd_sc_hd__nor2_8
XFILLER_109_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10370_ _11711_/CLK _10370_/D vssd1 vssd1 vccd1 vccd1 _10370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09029_ _11365_/Q _09035_/B vssd1 vssd1 vccd1 vccd1 _09029_/X sky130_fd_sc_hd__or2_1
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout750 _06589_/A2 vssd1 vssd1 vccd1 vccd1 _06504_/B1 sky130_fd_sc_hd__buf_4
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout761 _05749_/X vssd1 vssd1 vccd1 vccd1 _06674_/A2 sky130_fd_sc_hd__buf_6
Xfanout772 fanout782/X vssd1 vssd1 vccd1 vccd1 _07111_/A sky130_fd_sc_hd__buf_6
XFILLER_150_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout783 _07539_/A vssd1 vssd1 vccd1 vccd1 _06856_/A2 sky130_fd_sc_hd__buf_6
Xfanout794 _05746_/X vssd1 vssd1 vccd1 vccd1 _08971_/A sky130_fd_sc_hd__buf_12
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_110 _07153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _10134_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_132 _10023_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_143 _05449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _07052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_176 _09292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_187 _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _10021_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11755_/CLK _11755_/D vssd1 vssd1 vccd1 vccd1 _11755_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10706_ _11472_/CLK _10706_/D vssd1 vssd1 vccd1 vccd1 _10706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11686_ _11733_/CLK _11686_/D vssd1 vssd1 vccd1 vccd1 _11686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10637_ _10644_/CLK _10637_/D vssd1 vssd1 vccd1 vccd1 _10637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10568_ _11462_/CLK _10568_/D vssd1 vssd1 vccd1 vccd1 _10568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10499_ _10804_/CLK _10499_/D vssd1 vssd1 vccd1 vccd1 _10499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput5 io_in[9] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
X_06730_ _10711_/Q _07777_/A _06875_/A2 _10782_/Q _06726_/X vssd1 vssd1 vccd1 vccd1
+ _06730_/X sky130_fd_sc_hd__o221a_1
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06661_ input84/X _06655_/X _06660_/X _06576_/A vssd1 vssd1 vccd1 vccd1 _06661_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05612_ _05616_/A1 _11396_/Q _11393_/Q _11626_/Q _05611_/X vssd1 vssd1 vccd1 vccd1
+ _05615_/A sky130_fd_sc_hd__a221o_4
X_08400_ _09995_/A1 _11041_/Q _08414_/S vssd1 vssd1 vccd1 vccd1 _08401_/B sky130_fd_sc_hd__mux2_1
X_09380_ _09380_/A _10108_/B _10180_/C vssd1 vssd1 vccd1 vccd1 _09390_/S sky130_fd_sc_hd__or3_4
X_06592_ _10450_/Q _07222_/A _10009_/A _11219_/Q vssd1 vssd1 vccd1 vccd1 _06592_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_149_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08331_ _11006_/Q _08323_/Y _08324_/Y _07314_/X vssd1 vssd1 vccd1 vccd1 _11006_/D
+ sky130_fd_sc_hd__o22a_1
X_05543_ _05543_/A _05543_/B vssd1 vssd1 vccd1 vccd1 _05543_/Y sky130_fd_sc_hd__nor2_8
XFILLER_51_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08262_ _09995_/A1 _10963_/Q _08272_/S vssd1 vssd1 vccd1 vccd1 _08263_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05474_ _05474_/A _05474_/B _06950_/A vssd1 vssd1 vccd1 vccd1 _05475_/D sky130_fd_sc_hd__or3_4
XFILLER_123_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07213_ _07025_/A _07204_/B _07771_/B1 _10370_/Q vssd1 vssd1 vccd1 vccd1 _10370_/D
+ sky130_fd_sc_hd__a22o_1
X_08193_ _08193_/A _08193_/B vssd1 vssd1 vccd1 vccd1 _10931_/D sky130_fd_sc_hd__or2_1
XFILLER_118_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07144_ _10333_/Q _07145_/B _07188_/S _07143_/X vssd1 vssd1 vccd1 vccd1 _10333_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_69_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07075_ _10050_/A _07075_/B vssd1 vssd1 vccd1 vccd1 _10296_/D sky130_fd_sc_hd__or2_1
XFILLER_134_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06026_ _11373_/Q _06221_/A2 _09110_/A _11406_/Q _06025_/X vssd1 vssd1 vccd1 vccd1
+ _06026_/X sky130_fd_sc_hd__o221a_2
XFILLER_86_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07977_ _10812_/Q _07092_/A _07977_/S vssd1 vssd1 vccd1 vccd1 _07978_/B sky130_fd_sc_hd__mux2_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09716_ _10415_/Q _09871_/A2 _09886_/B1 _11439_/Q _09715_/X vssd1 vssd1 vccd1 vccd1
+ _09721_/B sky130_fd_sc_hd__a221o_1
X_06928_ _09256_/A1 _10206_/Q _06934_/S vssd1 vssd1 vccd1 vccd1 _10206_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09647_ _10324_/Q _09944_/B1 _09646_/X vssd1 vssd1 vccd1 vccd1 _09650_/C sky130_fd_sc_hd__a21o_1
X_06859_ _10377_/Q _07904_/A _06858_/X _06873_/D1 vssd1 vssd1 vccd1 vccd1 _06859_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09578_ _10508_/Q _09568_/B _09571_/D _10509_/Q vssd1 vssd1 vccd1 vccd1 _09578_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08789_/A1 _11114_/Q _08529_/S vssd1 vssd1 vccd1 vccd1 _08530_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ _11800_/CLK _11540_/D vssd1 vssd1 vccd1 vccd1 _11540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11471_ _11471_/CLK _11471_/D vssd1 vssd1 vccd1 vccd1 _11471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10422_ _10644_/CLK _10422_/D vssd1 vssd1 vccd1 vccd1 _10422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10353_ _10808_/CLK _10353_/D vssd1 vssd1 vccd1 vccd1 _10353_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_100_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10284_ _11698_/CLK _10284_/D vssd1 vssd1 vccd1 vccd1 _10284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout580 _05819_/Y vssd1 vssd1 vccd1 vccd1 _06665_/A2 sky130_fd_sc_hd__buf_2
Xfanout591 _09959_/A vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__buf_6
XFILLER_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _11808_/CLK _11807_/D vssd1 vssd1 vccd1 vccd1 _11807_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _11765_/CLK _11738_/D vssd1 vssd1 vccd1 vccd1 _11738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11669_ _11756_/CLK _11669_/D vssd1 vssd1 vccd1 vccd1 _11669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05190_ _05190_/A _05190_/B vssd1 vssd1 vccd1 vccd1 _05190_/Y sky130_fd_sc_hd__nor2_4
XFILLER_127_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07900_ _07039_/A _07966_/S _07899_/X _07902_/C1 vssd1 vssd1 vccd1 vccd1 _10768_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08880_ _08933_/A1 _11297_/Q _08890_/S vssd1 vssd1 vccd1 vccd1 _08881_/B sky130_fd_sc_hd__mux2_1
XFILLER_57_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07831_ _08661_/A _07820_/B _07821_/A _10726_/Q vssd1 vssd1 vccd1 vccd1 _10726_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07762_ _10682_/Q _08441_/B2 _07773_/S vssd1 vssd1 vccd1 vccd1 _10682_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09501_ _09501_/A vssd1 vssd1 vccd1 vccd1 _09501_/Y sky130_fd_sc_hd__inv_2
X_06713_ _10293_/Q _06873_/A2 _06685_/B _11713_/Q _06712_/X vssd1 vssd1 vccd1 vccd1
+ _06713_/X sky130_fd_sc_hd__o221a_1
X_07693_ _08655_/B _08591_/B vssd1 vssd1 vccd1 vccd1 _07693_/Y sky130_fd_sc_hd__nor2_2
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06644_ _07083_/A _06644_/B _06644_/C vssd1 vssd1 vccd1 vccd1 _06644_/X sky130_fd_sc_hd__or3_4
X_09432_ _09681_/B _09432_/B vssd1 vssd1 vccd1 vccd1 _09692_/B sky130_fd_sc_hd__or2_4
XFILLER_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09363_ _11539_/Q _09359_/X _09362_/X vssd1 vssd1 vccd1 vccd1 _11539_/D sky130_fd_sc_hd__a21o_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06575_ input85/X _06569_/X _06574_/X _11871_/A vssd1 vssd1 vccd1 vccd1 _06576_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05526_ _05616_/A1 _11505_/Q _11502_/Q _05077_/A vssd1 vssd1 vccd1 vccd1 _05526_/X
+ sky130_fd_sc_hd__a22o_1
X_08314_ _10111_/A0 _10993_/Q _08321_/S vssd1 vssd1 vccd1 vccd1 _10993_/D sky130_fd_sc_hd__mux2_1
X_09294_ _10161_/A1 _09310_/B _10166_/B1 vssd1 vssd1 vccd1 vccd1 _09294_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_10 _05734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_21 _06568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 _07022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ _08245_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08245_/X sky130_fd_sc_hd__or2_4
XANTENNA_54 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05457_ _10758_/Q _09881_/A2 _09878_/B1 _10759_/Q vssd1 vssd1 vccd1 vccd1 _05457_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_65 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_76 _11615_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_87 _08440_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08176_ _07057_/A _10918_/Q _08181_/S vssd1 vssd1 vccd1 vccd1 _10918_/D sky130_fd_sc_hd__mux2_1
XANTENNA_98 _09572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05388_ _10473_/Q _10472_/Q _05399_/S vssd1 vssd1 vccd1 vccd1 _05389_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_1324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07127_ _10134_/A0 _07111_/X _07126_/X _07107_/B vssd1 vssd1 vccd1 vccd1 _10323_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07058_ _10287_/Q _07047_/B _07490_/S _07314_/B vssd1 vssd1 vccd1 vccd1 _10287_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput150 _11573_/Q vssd1 vssd1 vccd1 vccd1 ram_addr[4] sky130_fd_sc_hd__buf_4
XFILLER_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput161 _11581_/Q vssd1 vssd1 vccd1 vccd1 rom_addr[3] sky130_fd_sc_hd__buf_4
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput172 _11870_/X vssd1 vssd1 vccd1 vccd1 wb_rom_adrb[4] sky130_fd_sc_hd__buf_4
X_06009_ _10592_/Q _06539_/B1 _06008_/X _06265_/C1 vssd1 vssd1 vccd1 vccd1 _06009_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput183 _05489_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_4
XFILLER_82_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput194 _05499_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_4
XFILLER_99_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10971_ _11575_/CLK _10971_/D vssd1 vssd1 vccd1 vccd1 _10971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11523_ _11685_/CLK _11523_/D vssd1 vssd1 vccd1 vccd1 _11523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11454_ _11661_/CLK _11454_/D vssd1 vssd1 vccd1 vccd1 _11454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10405_ _10666_/CLK _10405_/D vssd1 vssd1 vccd1 vccd1 _10405_/Q sky130_fd_sc_hd__dfxtp_1
X_11385_ _11385_/CLK _11385_/D vssd1 vssd1 vccd1 vccd1 _11385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10336_ _11474_/CLK _10336_/D vssd1 vssd1 vccd1 vccd1 _10336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _11698_/CLK _10267_/D vssd1 vssd1 vccd1 vccd1 _10267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10198_ _11810_/CLK _10198_/D vssd1 vssd1 vccd1 vccd1 _10198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_128_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10725_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06360_ _11547_/Q _09359_/A _06413_/A2 _11755_/Q vssd1 vssd1 vccd1 vccd1 _06360_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05311_ _11018_/Q _11017_/Q _05377_/S vssd1 vssd1 vccd1 vccd1 _05312_/D sky130_fd_sc_hd__mux2_1
X_06291_ _11347_/Q _08972_/A _06718_/B1 _11420_/Q vssd1 vssd1 vccd1 vccd1 _06291_/X
+ sky130_fd_sc_hd__o22a_1
X_08030_ _10178_/A1 _08027_/S _08029_/X _07011_/B vssd1 vssd1 vccd1 vccd1 _10839_/D
+ sky130_fd_sc_hd__o211a_1
X_05242_ _10794_/Q _10793_/Q _05419_/S vssd1 vssd1 vccd1 vccd1 _05248_/C sky130_fd_sc_hd__mux2_2
Xinput30 rom_value[28] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_2
Xinput41 rom_value[9] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput52 wb_rom_val[19] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_4
Xinput63 wb_rom_val[29] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_4
Xinput74 wb_rst_i vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_12
X_05173_ _11228_/Q _11227_/Q _05398_/S vssd1 vssd1 vccd1 vccd1 _05178_/C sky130_fd_sc_hd__mux2_1
Xinput85 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__buf_4
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput96 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09981_ _10162_/A1 _09977_/X _09980_/X _09995_/C1 vssd1 vssd1 vccd1 vccd1 _11677_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08932_ _11325_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08932_/X sky130_fd_sc_hd__or2_1
XFILLER_130_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08863_ _08873_/A _08863_/B vssd1 vssd1 vccd1 vccd1 _11288_/D sky130_fd_sc_hd__or2_1
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07814_ _07934_/A _07814_/B vssd1 vssd1 vccd1 vccd1 _10714_/D sky130_fd_sc_hd__or2_1
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08794_ _11253_/Q _08804_/B vssd1 vssd1 vccd1 vccd1 _08794_/X sky130_fd_sc_hd__or2_1
XFILLER_26_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07745_ _07932_/A1 _07761_/A2 _07744_/X _07932_/C1 vssd1 vssd1 vccd1 vccd1 _10673_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07676_ _08438_/A _08663_/S vssd1 vssd1 vccd1 vccd1 _07676_/X sky130_fd_sc_hd__or2_4
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09415_ _11604_/Q _11603_/Q vssd1 vssd1 vccd1 vccd1 _09416_/B sky130_fd_sc_hd__nor2_2
X_06627_ _11032_/Q _10087_/A _06623_/X _06626_/X vssd1 vssd1 vccd1 vccd1 _06633_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ _11527_/Q _09326_/X _09345_/X vssd1 vssd1 vccd1 vccd1 _11527_/D sky130_fd_sc_hd__a21o_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06558_ _06554_/X _06557_/X _06431_/A _06552_/X vssd1 vssd1 vccd1 vccd1 _06558_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_40_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05509_ input2/X _11335_/Q _10213_/Q vssd1 vssd1 vccd1 vccd1 _11605_/D sky130_fd_sc_hd__mux2_1
X_09277_ _11490_/Q _09271_/X _09276_/X vssd1 vssd1 vccd1 vccd1 _11490_/D sky130_fd_sc_hd__a21o_1
X_06489_ _11114_/Q _06646_/A2 _06487_/X _06488_/X vssd1 vssd1 vccd1 vccd1 _06489_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08228_ _08469_/A _08225_/S _08227_/X _08351_/C1 vssd1 vssd1 vccd1 vccd1 _10948_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08159_ _08757_/A _08159_/B vssd1 vssd1 vccd1 vccd1 _10905_/D sky130_fd_sc_hd__or2_1
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11170_ _11325_/CLK _11170_/D vssd1 vssd1 vccd1 vccd1 _11170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10121_ _07002_/A _11767_/Q _10135_/S vssd1 vssd1 vccd1 vccd1 _11767_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10052_ _10058_/A _10052_/B vssd1 vssd1 vccd1 vccd1 _11717_/D sky130_fd_sc_hd__or2_1
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10954_ _11485_/CLK _10954_/D vssd1 vssd1 vccd1 vccd1 _10954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10885_ _10932_/CLK _10885_/D vssd1 vssd1 vccd1 vccd1 _10885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11506_ _11800_/CLK _11506_/D vssd1 vssd1 vccd1 vccd1 _11506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11437_ _11458_/CLK _11437_/D vssd1 vssd1 vccd1 vccd1 _11437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11368_ _11808_/CLK _11368_/D vssd1 vssd1 vccd1 vccd1 _11368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _11710_/CLK _10319_/D vssd1 vssd1 vccd1 vccd1 _10319_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _11332_/CLK _11299_/D vssd1 vssd1 vccd1 vccd1 _11299_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05860_ _10617_/Q _06371_/A2 _07827_/A2 _10976_/Q vssd1 vssd1 vccd1 vccd1 _05860_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05791_ _11313_/Q _09271_/A _06716_/B1 _11239_/Q _05790_/X vssd1 vssd1 vccd1 vccd1
+ _05791_/X sky130_fd_sc_hd__o221a_1
XFILLER_19_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07530_ _07918_/A _07530_/B vssd1 vssd1 vccd1 vccd1 _10549_/D sky130_fd_sc_hd__or2_1
XFILLER_81_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07461_ _10017_/A0 _10508_/Q _07477_/S vssd1 vssd1 vccd1 vccd1 _07462_/B sky130_fd_sc_hd__mux2_1
XFILLER_74_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09200_ input106/X _11447_/Q _09200_/S vssd1 vssd1 vccd1 vccd1 _09200_/X sky130_fd_sc_hd__mux2_1
X_06412_ _10589_/Q _06454_/A2 _06412_/B1 _10840_/Q _06624_/C1 vssd1 vssd1 vccd1 vccd1
+ _06412_/X sky130_fd_sc_hd__o221a_1
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07392_ _08193_/A _07392_/B vssd1 vssd1 vccd1 vccd1 _10472_/D sky130_fd_sc_hd__or2_1
XFILLER_148_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09131_ _09131_/A _10136_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09149_/B sky130_fd_sc_hd__and3_4
X_06343_ _11675_/Q _09965_/A _09380_/A _11000_/Q vssd1 vssd1 vccd1 vccd1 _06343_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09062_ _11379_/Q _09060_/X _09061_/X vssd1 vssd1 vccd1 vccd1 _11379_/D sky130_fd_sc_hd__a21o_1
XFILLER_124_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06274_ _07082_/A _06272_/X _06273_/X _05816_/A vssd1 vssd1 vccd1 vccd1 _06274_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_96_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11442_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08013_ _10831_/Q _08091_/C vssd1 vssd1 vccd1 vccd1 _08013_/X sky130_fd_sc_hd__or2_1
X_05225_ _05413_/S _11007_/Q vssd1 vssd1 vccd1 vccd1 _05225_/X sky130_fd_sc_hd__and2_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11634_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05156_ _05156_/A _05156_/B _05156_/C _05156_/D vssd1 vssd1 vccd1 vccd1 _05157_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_143_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09964_ _09827_/Y _09963_/B _09963_/Y vssd1 vssd1 vccd1 vccd1 _11665_/D sky130_fd_sc_hd__a21oi_1
X_05087_ _06939_/A vssd1 vssd1 vccd1 vccd1 _09539_/A sky130_fd_sc_hd__inv_6
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08915_ _09090_/A1 _08945_/A2 _08914_/X _09078_/C1 vssd1 vssd1 vccd1 vccd1 _11316_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _11744_/Q _09566_/D _09573_/D _11701_/Q vssd1 vssd1 vccd1 vccd1 _09895_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _08846_/A0 _11281_/Q _08850_/S vssd1 vssd1 vccd1 vccd1 _08847_/B sky130_fd_sc_hd__mux2_1
XFILLER_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _09283_/A1 _08802_/S _08776_/X _08919_/C1 vssd1 vssd1 vccd1 vccd1 _11244_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_73_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05989_ _11192_/Q _06736_/A2 _06735_/B1 _11155_/Q _05988_/X vssd1 vssd1 vccd1 vccd1
+ _05989_/X sky130_fd_sc_hd__o221a_2
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _10665_/Q _07760_/B vssd1 vssd1 vccd1 vccd1 _07728_/X sky130_fd_sc_hd__or2_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07659_ _07659_/A _07659_/B vssd1 vssd1 vccd1 vccd1 _10622_/D sky130_fd_sc_hd__or2_1
XFILLER_43_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10670_ _10773_/CLK _10670_/D vssd1 vssd1 vccd1 vccd1 _10670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09329_ _11519_/Q _09343_/B vssd1 vssd1 vccd1 vccd1 _09329_/X sky130_fd_sc_hd__or2_1
XFILLER_16_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11222_ _11629_/CLK _11222_/D vssd1 vssd1 vccd1 vccd1 _11222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ _11393_/CLK _11153_/D vssd1 vssd1 vccd1 vccd1 _11153_/Q sky130_fd_sc_hd__dfxtp_1
X_10104_ _11754_/Q _10104_/B vssd1 vssd1 vccd1 vccd1 _10104_/X sky130_fd_sc_hd__or2_1
XFILLER_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11084_ _11140_/CLK _11084_/D vssd1 vssd1 vccd1 vccd1 _11084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10035_ _10039_/A _10035_/B vssd1 vssd1 vccd1 vccd1 _11707_/D sky130_fd_sc_hd__or2_1
XFILLER_88_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10937_ _11312_/CLK _10937_/D vssd1 vssd1 vccd1 vccd1 _10937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10868_ _11485_/CLK _10868_/D vssd1 vssd1 vccd1 vccd1 _10868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10799_ _11477_/CLK _10799_/D vssd1 vssd1 vccd1 vccd1 _10799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout409 _05379_/Y vssd1 vssd1 vccd1 vccd1 _09565_/C sky130_fd_sc_hd__buf_4
XFILLER_63_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06961_ _11607_/Q _09538_/C _06944_/A _09488_/C vssd1 vssd1 vccd1 vccd1 _06961_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08700_ _08853_/A1 _08695_/S _08699_/X _08937_/C1 vssd1 vssd1 vccd1 vccd1 _11204_/D
+ sky130_fd_sc_hd__o211a_1
X_05912_ _10523_/Q _06106_/B _05908_/X _05911_/X vssd1 vssd1 vccd1 vccd1 _05912_/X
+ sky130_fd_sc_hd__o211a_1
X_09680_ _11604_/Q _09680_/B _09680_/C _11603_/Q vssd1 vssd1 vccd1 vccd1 _09681_/D
+ sky130_fd_sc_hd__or4b_1
X_06892_ _06892_/A _06892_/B vssd1 vssd1 vccd1 vccd1 _08243_/C sky130_fd_sc_hd__or2_4
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_143_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11779_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08631_ _11170_/Q _08633_/B vssd1 vssd1 vccd1 vccd1 _08631_/X sky130_fd_sc_hd__or2_1
X_05843_ _07690_/A _05842_/X _05832_/X _05095_/Y vssd1 vssd1 vccd1 vccd1 _05843_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08562_ _08733_/A _08562_/B vssd1 vssd1 vccd1 vccd1 _11135_/D sky130_fd_sc_hd__or2_1
XFILLER_78_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05774_ _08243_/A _11872_/A vssd1 vssd1 vccd1 vccd1 _05774_/Y sky130_fd_sc_hd__nor2_4
XFILLER_39_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07513_ _08846_/A0 _10541_/Q _07513_/S vssd1 vssd1 vccd1 vccd1 _07514_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08493_ _11097_/Q _08503_/B vssd1 vssd1 vccd1 vccd1 _08493_/X sky130_fd_sc_hd__or2_1
XFILLER_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07444_ _10496_/Q _07441_/Y _07443_/Y _08440_/B2 vssd1 vssd1 vccd1 vccd1 _10496_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07375_ _08050_/A _07393_/S vssd1 vssd1 vccd1 vccd1 _07655_/S sky130_fd_sc_hd__nor2_8
XFILLER_149_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09114_ _09114_/A1 _09110_/X _09113_/X _09279_/C1 vssd1 vssd1 vccd1 vccd1 _11403_/D
+ sky130_fd_sc_hd__o211a_1
X_06326_ _11095_/Q _06629_/B1 _06325_/X _06392_/C1 vssd1 vssd1 vccd1 vccd1 _06326_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09045_ _11372_/Q _09055_/B vssd1 vssd1 vccd1 vccd1 _09045_/X sky130_fd_sc_hd__or2_1
XFILLER_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06257_ _10916_/Q _08166_/A _06636_/A2 _11076_/Q _06256_/X vssd1 vssd1 vccd1 vccd1
+ _06257_/X sky130_fd_sc_hd__o221a_1
X_05208_ _10434_/Q _10433_/Q _05419_/S vssd1 vssd1 vccd1 vccd1 _05214_/C sky130_fd_sc_hd__mux2_2
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06188_ _10209_/Q _06351_/A2 _06184_/X _06187_/X vssd1 vssd1 vccd1 vccd1 _06188_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05139_ _10638_/Q _10637_/Q _05416_/S vssd1 vssd1 vccd1 vccd1 _05140_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout910 _05093_/Y vssd1 vssd1 vccd1 vccd1 _06577_/A sky130_fd_sc_hd__buf_6
XFILLER_85_1299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout921 _06297_/C1 vssd1 vssd1 vccd1 vccd1 _06624_/C1 sky130_fd_sc_hd__clkbuf_8
Xfanout932 _10162_/A1 vssd1 vssd1 vccd1 vccd1 _09114_/A1 sky130_fd_sc_hd__buf_4
X_09947_ _10367_/Q _09947_/A2 _09947_/B1 _10693_/Q vssd1 vssd1 vccd1 vccd1 _09947_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout943 input95/X vssd1 vssd1 vccd1 vccd1 _09216_/A0 sky130_fd_sc_hd__clkbuf_16
Xfanout954 fanout958/X vssd1 vssd1 vccd1 vccd1 _08760_/A0 sky130_fd_sc_hd__buf_2
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout965 _08933_/A1 vssd1 vssd1 vccd1 vccd1 _07104_/A sky130_fd_sc_hd__buf_12
XFILLER_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout976 _10181_/A0 vssd1 vssd1 vccd1 vccd1 _09999_/A0 sky130_fd_sc_hd__buf_6
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _10575_/Q _09878_/A2 _09878_/B1 _10571_/Q vssd1 vssd1 vccd1 vccd1 _09878_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout987 _11870_/A vssd1 vssd1 vccd1 vccd1 _07689_/A sky130_fd_sc_hd__buf_12
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout998 _06670_/D1 vssd1 vssd1 vccd1 vccd1 _06873_/D1 sky130_fd_sc_hd__buf_8
XFILLER_85_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08829_ _10190_/A0 _08838_/S _08828_/X _08841_/C1 vssd1 vssd1 vccd1 vccd1 _11272_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11780_/CLK _11771_/D vssd1 vssd1 vccd1 vccd1 _11771_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1089 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1089/HI io_oeb[19] sky130_fd_sc_hd__conb_1
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10722_ _10798_/CLK _10722_/D vssd1 vssd1 vccd1 vccd1 _10722_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653_ _11067_/CLK _10653_/D vssd1 vssd1 vccd1 vccd1 _10653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10584_ _11628_/CLK _10584_/D vssd1 vssd1 vccd1 vccd1 _10584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11205_ _11329_/CLK _11205_/D vssd1 vssd1 vccd1 vccd1 _11205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11136_ _11136_/CLK _11136_/D vssd1 vssd1 vccd1 vccd1 _11136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11067_ _11067_/CLK _11067_/D vssd1 vssd1 vccd1 vccd1 _11067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10018_ _10020_/A _10018_/B vssd1 vssd1 vccd1 vccd1 _11699_/D sky130_fd_sc_hd__or2_1
XFILLER_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05490_ _10235_/Q input46/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05490_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07160_ _07785_/A0 _10341_/Q _09243_/C vssd1 vssd1 vccd1 vccd1 _07161_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06111_ _10399_/Q _06804_/B _07455_/A _10658_/Q vssd1 vssd1 vccd1 vccd1 _06111_/X
+ sky130_fd_sc_hd__o22a_1
X_07091_ _10301_/Q _07090_/X _07109_/S vssd1 vssd1 vccd1 vccd1 _10301_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06042_ _10524_/Q _06308_/A2 _06373_/B1 _10314_/Q _06041_/X vssd1 vssd1 vccd1 vccd1
+ _06042_/X sky130_fd_sc_hd__o221a_2
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout217 _07624_/Y vssd1 vssd1 vccd1 vccd1 _07626_/S sky130_fd_sc_hd__buf_2
X_09801_ _10523_/Q _09566_/B _09571_/D _10283_/Q vssd1 vssd1 vccd1 vccd1 _09801_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout228 _07188_/S vssd1 vssd1 vccd1 vccd1 _07186_/S sky130_fd_sc_hd__buf_6
XFILLER_59_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout239 _10009_/Y vssd1 vssd1 vccd1 vccd1 _10057_/S sky130_fd_sc_hd__clkbuf_4
X_07993_ _09325_/A _08649_/C _09037_/C vssd1 vssd1 vccd1 vccd1 _08091_/C sky130_fd_sc_hd__and3_4
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09732_ _11474_/Q _09879_/A2 _09567_/D _10348_/Q vssd1 vssd1 vccd1 vccd1 _09732_/X
+ sky130_fd_sc_hd__a22o_1
X_06944_ _06944_/A vssd1 vssd1 vccd1 vccd1 _06944_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09663_ _09599_/X _09618_/X _09640_/X _09959_/B vssd1 vssd1 vccd1 vccd1 _09665_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06875_ _11463_/Q _06875_/A2 _06875_/B1 _10681_/Q vssd1 vssd1 vccd1 vccd1 _06875_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08614_ _08682_/A _08614_/B vssd1 vssd1 vccd1 vccd1 _11161_/D sky130_fd_sc_hd__or2_1
X_05826_ _11793_/Q _10159_/A _09977_/A _11677_/Q _05825_/X vssd1 vssd1 vccd1 vccd1
+ _05826_/X sky130_fd_sc_hd__o221a_1
XFILLER_27_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09594_ _11658_/Q _09594_/B _09594_/C _09594_/D vssd1 vssd1 vccd1 vccd1 _09594_/X
+ sky130_fd_sc_hd__and4_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08545_ _11122_/Q _08545_/B vssd1 vssd1 vccd1 vccd1 _08545_/X sky130_fd_sc_hd__or2_1
X_05757_ _11389_/Q _06219_/A2 _09132_/A _11412_/Q vssd1 vssd1 vccd1 vccd1 _05757_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08476_ _09393_/A0 _08497_/S _08475_/X _09022_/C1 vssd1 vssd1 vccd1 vccd1 _11088_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05688_ _11161_/Q _05573_/Y _05579_/Y _11168_/Q _05687_/X vssd1 vssd1 vccd1 vccd1
+ _05691_/B sky130_fd_sc_hd__a221o_2
XFILLER_23_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07427_ _10047_/A1 _10490_/Q _07437_/S vssd1 vssd1 vccd1 vccd1 _07428_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11675_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_136_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07358_ _09248_/A _08649_/B _08560_/C vssd1 vssd1 vccd1 vccd1 _07977_/S sky130_fd_sc_hd__and3_4
XFILLER_109_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06309_ _06309_/A _06309_/B _06309_/C vssd1 vssd1 vccd1 vccd1 _06309_/X sky130_fd_sc_hd__and3_2
XFILLER_136_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07289_ _07141_/A _10413_/Q _09184_/S vssd1 vssd1 vccd1 vccd1 _07290_/B sky130_fd_sc_hd__mux2_1
XFILLER_124_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09028_ _10149_/A1 _09016_/X _09027_/X _09036_/C1 vssd1 vssd1 vccd1 vccd1 _11364_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout740 _09292_/A vssd1 vssd1 vccd1 vccd1 _09109_/A sky130_fd_sc_hd__buf_8
XFILLER_49_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout751 _06214_/B1 vssd1 vssd1 vccd1 vccd1 _06589_/A2 sky130_fd_sc_hd__buf_6
Xfanout762 _06718_/B1 vssd1 vssd1 vccd1 vccd1 _08855_/A sky130_fd_sc_hd__buf_6
Xfanout773 fanout782/X vssd1 vssd1 vccd1 vccd1 _06373_/B1 sky130_fd_sc_hd__buf_4
Xfanout784 fanout793/X vssd1 vssd1 vccd1 vccd1 _07539_/A sky130_fd_sc_hd__buf_6
XFILLER_74_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout795 _05746_/X vssd1 vssd1 vccd1 vccd1 _09248_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_92_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_100 _09566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _09976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 fanout958/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_133 _10019_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_144 _05730_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_155 _07105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _06674_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11791_/CLK _11754_/D vssd1 vssd1 vccd1 vccd1 _11754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_188 _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _10021_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _10765_/CLK _10705_/D vssd1 vssd1 vccd1 vccd1 _10705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11685_ _11685_/CLK _11685_/D vssd1 vssd1 vccd1 vccd1 _11685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10636_ _10644_/CLK _10636_/D vssd1 vssd1 vccd1 vccd1 _10636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10567_ _11575_/CLK _10567_/D vssd1 vssd1 vccd1 vccd1 _10567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10498_ _10804_/CLK _10498_/D vssd1 vssd1 vccd1 vccd1 _10498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11119_ _11572_/CLK _11119_/D vssd1 vssd1 vccd1 vccd1 _11119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput6 ram_val_in[0] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_4
XFILLER_77_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06660_ _11167_/Q _09037_/A _06656_/X _06659_/X vssd1 vssd1 vccd1 vccd1 _06660_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05611_ _05618_/A1 _11392_/Q _11389_/Q _11624_/Q vssd1 vssd1 vccd1 vccd1 _05611_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06591_ _10923_/Q _06591_/A2 _06635_/B1 _11267_/Q vssd1 vssd1 vccd1 vccd1 _06591_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_64_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08330_ _11005_/Q _08322_/Y _08325_/Y _09232_/B2 vssd1 vssd1 vccd1 vccd1 _11005_/D
+ sky130_fd_sc_hd__a22o_1
X_05542_ _05626_/A2 _11355_/Q _11350_/Q _05630_/B1 _05541_/X vssd1 vssd1 vccd1 vccd1
+ _05543_/B sky130_fd_sc_hd__a221o_4
XFILLER_75_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05473_ _09538_/A _05473_/B vssd1 vssd1 vccd1 vccd1 _06950_/A sky130_fd_sc_hd__nor2_2
X_08261_ _08987_/A1 _08276_/S _08260_/X _08921_/C1 vssd1 vssd1 vccd1 vccd1 _10962_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07212_ _07211_/A _07205_/B _07773_/S _10369_/Q vssd1 vssd1 vccd1 vccd1 _10369_/D
+ sky130_fd_sc_hd__o22a_1
X_08192_ _10931_/Q _10132_/A0 _08197_/S vssd1 vssd1 vccd1 vccd1 _08193_/B sky130_fd_sc_hd__mux2_1
X_07143_ _07143_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _07143_/X sky130_fd_sc_hd__and2_4
XFILLER_106_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07074_ _07034_/A _10296_/Q _07074_/S vssd1 vssd1 vccd1 vccd1 _07075_/B sky130_fd_sc_hd__mux2_1
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06025_ _11492_/Q _09271_/A _08972_/A _11343_/Q vssd1 vssd1 vccd1 vccd1 _06025_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07976_ _08733_/A _07976_/B vssd1 vssd1 vccd1 vccd1 _10811_/D sky130_fd_sc_hd__or2_1
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09715_ _10409_/Q _09883_/B1 _09565_/C _11436_/Q _09714_/X vssd1 vssd1 vccd1 vccd1
+ _09715_/X sky130_fd_sc_hd__a221o_1
XFILLER_68_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06927_ _10111_/A0 _10205_/Q _06934_/S vssd1 vssd1 vccd1 vccd1 _10205_/D sky130_fd_sc_hd__mux2_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09646_ _10334_/Q _09567_/A _09573_/B _10319_/Q vssd1 vssd1 vccd1 vccd1 _09646_/X
+ sky130_fd_sc_hd__a22o_1
X_06858_ _10299_/Q _06873_/A2 _06858_/B1 _10278_/Q _06857_/X vssd1 vssd1 vccd1 vccd1
+ _06858_/X sky130_fd_sc_hd__o221a_1
XFILLER_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05809_ _11053_/Q _08054_/A _08123_/A _10888_/Q _06392_/C1 vssd1 vssd1 vccd1 vccd1
+ _05809_/X sky130_fd_sc_hd__o221a_1
XFILLER_93_1310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _10278_/Q _09568_/A _09953_/B1 _10279_/Q vssd1 vssd1 vccd1 vccd1 _09577_/X
+ sky130_fd_sc_hd__a22o_1
X_06789_ _10628_/Q _06871_/A2 _06785_/X _06788_/X vssd1 vssd1 vccd1 vccd1 _06789_/X
+ sky130_fd_sc_hd__o211a_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08528_ _08682_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _11113_/D sky130_fd_sc_hd__or2_1
XFILLER_93_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08459_ _11080_/Q _10135_/A0 _08459_/S vssd1 vssd1 vccd1 vccd1 _08460_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11470_ _11470_/CLK _11470_/D vssd1 vssd1 vccd1 vccd1 _11470_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_104_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10421_ _11233_/CLK _10421_/D vssd1 vssd1 vccd1 vccd1 _10421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10352_ _10769_/CLK _10352_/D vssd1 vssd1 vccd1 vccd1 _10352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10283_ _11703_/CLK _10283_/D vssd1 vssd1 vccd1 vccd1 _10283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout570 _08682_/A vssd1 vssd1 vccd1 vccd1 _08875_/A sky130_fd_sc_hd__clkbuf_4
Xfanout581 _05819_/Y vssd1 vssd1 vccd1 vccd1 _06704_/B sky130_fd_sc_hd__buf_6
XFILLER_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout592 _05101_/Y vssd1 vssd1 vccd1 vccd1 _09959_/A sky130_fd_sc_hd__buf_12
XFILLER_150_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _11808_/CLK _11806_/D vssd1 vssd1 vccd1 vccd1 _11806_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11762_/CLK _11737_/D vssd1 vssd1 vccd1 vccd1 _11737_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11668_ _11758_/CLK _11668_/D vssd1 vssd1 vccd1 vccd1 _11668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10619_ _11310_/CLK _10619_/D vssd1 vssd1 vccd1 vccd1 _10619_/Q sky130_fd_sc_hd__dfxtp_1
X_11599_ _11601_/CLK _11599_/D vssd1 vssd1 vccd1 vccd1 _11599_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07830_ _07104_/A _07820_/B _07821_/A _10725_/Q vssd1 vssd1 vccd1 vccd1 _10725_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07761_ _07042_/A _07761_/A2 _07760_/X _07932_/C1 vssd1 vssd1 vccd1 vccd1 _10681_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09500_ _09528_/A _09500_/B _09500_/C vssd1 vssd1 vccd1 vccd1 _09501_/A sky130_fd_sc_hd__nand3_1
XFILLER_38_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06712_ _10371_/Q _07203_/A _06872_/A2 _10489_/Q vssd1 vssd1 vccd1 vccd1 _06712_/X
+ sky130_fd_sc_hd__o22a_1
X_07692_ _07692_/A _08665_/C _09038_/C vssd1 vssd1 vccd1 vccd1 _08589_/S sky130_fd_sc_hd__or3_4
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09431_ _09477_/A _09431_/B _09554_/B _09672_/B vssd1 vssd1 vccd1 vccd1 _09432_/B
+ sky130_fd_sc_hd__or4_1
X_06643_ _10852_/Q _06643_/A2 _06639_/X _06642_/X vssd1 vssd1 vccd1 vccd1 _06644_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09362_ _10162_/A1 _09376_/B _10178_/B1 vssd1 vssd1 vccd1 vccd1 _09362_/X sky130_fd_sc_hd__a21o_1
XFILLER_75_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06574_ _11165_/Q _06649_/A2 _06570_/X _06573_/X vssd1 vssd1 vccd1 vccd1 _06574_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_33_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08313_ _10110_/A0 _10992_/Q _08321_/S vssd1 vssd1 vccd1 vccd1 _10992_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05525_ _11332_/Q _05518_/Y _05524_/Y _11323_/Q vssd1 vssd1 vccd1 vccd1 _05525_/X
+ sky130_fd_sc_hd__a22o_1
X_09293_ _09293_/A _10137_/B _10159_/C vssd1 vssd1 vccd1 vccd1 _09293_/X sky130_fd_sc_hd__or3_4
XFILLER_127_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_11 _05736_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_22 _06644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 _07303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ _08972_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08284_/B sky130_fd_sc_hd__nor2_8
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_44 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05456_ _10748_/Q _09875_/A2 _09875_/B1 _10747_/Q _05453_/X vssd1 vssd1 vccd1 vccd1
+ _05469_/B sky130_fd_sc_hd__a221o_1
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_55 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_66 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_77 _11615_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _10128_/A0 _10917_/Q _08181_/S vssd1 vssd1 vccd1 vccd1 _10917_/D sky130_fd_sc_hd__mux2_1
XANTENNA_88 _08440_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05387_ _10463_/Q _10462_/Q _05396_/S vssd1 vssd1 vccd1 vccd1 _05389_/C sky130_fd_sc_hd__mux2_1
XANTENNA_99 _09568_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ _10323_/Q _07126_/B vssd1 vssd1 vccd1 vccd1 _07126_/X sky130_fd_sc_hd__or2_1
XFILLER_106_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07057_ _07057_/A _07107_/B vssd1 vssd1 vccd1 vccd1 _07057_/X sky130_fd_sc_hd__and2_2
Xoutput140 _11620_/Q vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__buf_4
Xoutput151 _11574_/Q vssd1 vssd1 vccd1 vccd1 ram_addr[5] sky130_fd_sc_hd__buf_4
XFILLER_133_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput162 _11582_/Q vssd1 vssd1 vccd1 vccd1 rom_addr[4] sky130_fd_sc_hd__buf_4
X_06008_ _11234_/Q _06541_/A2 _06540_/A2 _10788_/Q _06007_/X vssd1 vssd1 vccd1 vccd1
+ _06008_/X sky130_fd_sc_hd__o221a_1
XFILLER_134_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput173 _11871_/X vssd1 vssd1 vccd1 vccd1 wb_rom_adrb[5] sky130_fd_sc_hd__buf_4
XFILLER_102_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput184 _05490_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_4
XFILLER_114_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput195 _05500_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_4
XFILLER_87_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07959_ _07187_/X _10801_/Q _07959_/S vssd1 vssd1 vccd1 vccd1 _10801_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10970_ _11622_/CLK _10970_/D vssd1 vssd1 vccd1 vccd1 _10970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09629_ _10803_/Q _09909_/A2 _09573_/C _10732_/Q _09622_/X vssd1 vssd1 vccd1 vccd1
+ _09633_/A sky130_fd_sc_hd__a221o_1
XFILLER_28_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _11683_/CLK _11522_/D vssd1 vssd1 vccd1 vccd1 _11522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11453_ _11465_/CLK _11453_/D vssd1 vssd1 vccd1 vccd1 _11453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10404_ _11644_/CLK _10404_/D vssd1 vssd1 vccd1 vccd1 _10404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11384_ _11428_/CLK _11384_/D vssd1 vssd1 vccd1 vccd1 _11384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10335_ _11744_/CLK _10335_/D vssd1 vssd1 vccd1 vccd1 _10335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10266_ _11698_/CLK _10266_/D vssd1 vssd1 vccd1 vccd1 _10266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10197_ _11803_/CLK _10197_/D vssd1 vssd1 vccd1 vccd1 _10197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05310_ _11024_/Q _11023_/Q _09680_/B vssd1 vssd1 vccd1 vccd1 _05312_/C sky130_fd_sc_hd__mux2_1
X_06290_ _11397_/Q _09082_/A _09110_/A _11410_/Q vssd1 vssd1 vccd1 vccd1 _06290_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput20 rom_value[19] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_2
X_05241_ _10866_/Q _10865_/Q _05413_/S vssd1 vssd1 vccd1 vccd1 _05248_/B sky130_fd_sc_hd__mux2_2
Xinput31 rom_value[29] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput42 wb_rom_val[0] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_2
Xinput53 wb_rom_val[1] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_2
XFILLER_122_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput64 wb_rom_val[2] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_2
X_05172_ _11232_/Q _11231_/Q _09680_/B vssd1 vssd1 vccd1 vccd1 _05178_/B sky130_fd_sc_hd__mux2_2
XFILLER_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput75 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_4
Xinput86 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput97 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__buf_6
X_09980_ _11677_/Q _09994_/B vssd1 vssd1 vccd1 vccd1 _09980_/X sky130_fd_sc_hd__or2_1
XFILLER_118_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08931_ _08931_/A1 _08940_/S _08930_/X _09078_/C1 vssd1 vssd1 vccd1 vccd1 _11324_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08862_ _09090_/A1 _11288_/Q _08890_/S vssd1 vssd1 vccd1 vccd1 _08863_/B sky130_fd_sc_hd__mux2_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07813_ _07933_/A0 _10714_/Q _09193_/B vssd1 vssd1 vccd1 vccd1 _07814_/B sky130_fd_sc_hd__mux2_1
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08793_ _08793_/A _08793_/B vssd1 vssd1 vccd1 vccd1 _11252_/D sky130_fd_sc_hd__or2_1
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07744_ _10673_/Q _07760_/B vssd1 vssd1 vccd1 vccd1 _07744_/X sky130_fd_sc_hd__or2_1
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07675_ _08303_/A _08663_/S vssd1 vssd1 vccd1 vccd1 _07675_/Y sky130_fd_sc_hd__nor2_2
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09414_ _11657_/Q _11575_/Q _09414_/S vssd1 vssd1 vccd1 vccd1 _11575_/D sky130_fd_sc_hd__mux2_1
X_06626_ _10954_/Q _10137_/A _06624_/X _06625_/X vssd1 vssd1 vccd1 vccd1 _06626_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09345_ _10178_/A1 _09343_/B _08851_/A vssd1 vssd1 vccd1 vccd1 _09345_/X sky130_fd_sc_hd__a21o_1
X_06557_ _10471_/Q _06642_/A2 _06556_/X _06642_/C1 vssd1 vssd1 vccd1 vccd1 _06557_/X
+ sky130_fd_sc_hd__o211a_1
X_05508_ _10253_/Q input66/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05508_/X sky130_fd_sc_hd__mux2_2
X_09276_ _09276_/A1 _09288_/B _09290_/B1 vssd1 vssd1 vccd1 vccd1 _09276_/X sky130_fd_sc_hd__a21o_1
X_06488_ _11200_/Q _06645_/A2 _09292_/A _11250_/Q vssd1 vssd1 vccd1 vccd1 _06488_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08227_ _10948_/Q _08902_/C vssd1 vssd1 vccd1 vccd1 _08227_/X sky130_fd_sc_hd__or2_1
X_05439_ _10669_/Q _09565_/A _09570_/B _10670_/Q vssd1 vssd1 vccd1 vccd1 _05439_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08158_ _09995_/A1 _10905_/Q _08162_/S vssd1 vssd1 vccd1 vccd1 _08159_/B sky130_fd_sc_hd__mux2_1
XFILLER_88_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07109_ _10309_/Q _07108_/X _07109_/S vssd1 vssd1 vccd1 vccd1 _10309_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08089_ _10870_/Q _08437_/A _08011_/S _08303_/A vssd1 vssd1 vccd1 vccd1 _08089_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_107_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10120_ _07048_/A _11766_/Q _10134_/S vssd1 vssd1 vccd1 vccd1 _11766_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10051_ _11717_/Q _10051_/A1 _10051_/S vssd1 vssd1 vccd1 vccd1 _10052_/B sky130_fd_sc_hd__mux2_1
XFILLER_103_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10953_ _11485_/CLK _10953_/D vssd1 vssd1 vccd1 vccd1 _10953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10884_ _10929_/CLK _10884_/D vssd1 vssd1 vccd1 vccd1 _10884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ _11801_/CLK _11505_/D vssd1 vssd1 vccd1 vccd1 _11505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11436_ _11457_/CLK _11436_/D vssd1 vssd1 vccd1 vccd1 _11436_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11367_ _11811_/CLK _11367_/D vssd1 vssd1 vccd1 vccd1 _11367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10318_ _10812_/CLK _10318_/D vssd1 vssd1 vccd1 vccd1 _10318_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _11330_/CLK _11298_/D vssd1 vssd1 vccd1 vccd1 _11298_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ _11474_/CLK _10249_/D vssd1 vssd1 vccd1 vccd1 _10249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05790_ _10955_/Q _08972_/A _06718_/B1 _11285_/Q vssd1 vssd1 vccd1 vccd1 _05790_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07460_ _10507_/Q _07000_/B _07000_/Y _07324_/B vssd1 vssd1 vccd1 vccd1 _10507_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06411_ _10865_/Q _06455_/A2 _06455_/B1 _10431_/Q vssd1 vssd1 vccd1 vccd1 _06411_/X
+ sky130_fd_sc_hd__o22a_1
X_07391_ _10472_/Q _08818_/A1 _07393_/S vssd1 vssd1 vccd1 vccd1 _07392_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09130_ _11411_/Q _09110_/X _09129_/X vssd1 vssd1 vccd1 vccd1 _11411_/D sky130_fd_sc_hd__a21o_1
XFILLER_37_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06342_ _11812_/Q _06883_/B _06341_/X vssd1 vssd1 vccd1 vccd1 _10230_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09061_ _10161_/A1 _09077_/B _08771_/A vssd1 vssd1 vccd1 vccd1 _09061_/X sky130_fd_sc_hd__a21o_1
X_06273_ _06633_/A _06266_/X _06271_/X _06619_/A1 _06261_/X vssd1 vssd1 vccd1 vccd1
+ _06273_/X sky130_fd_sc_hd__o311a_1
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ _08835_/A _08012_/B vssd1 vssd1 vccd1 vccd1 _10830_/D sky130_fd_sc_hd__or2_1
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05224_ _05224_/A _05224_/B _05224_/C _05224_/D vssd1 vssd1 vccd1 vccd1 _05224_/Y
+ sky130_fd_sc_hd__nor4_4
XFILLER_50_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05155_ _10942_/Q _10941_/Q _05377_/S vssd1 vssd1 vccd1 vccd1 _05156_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09963_ _11665_/Q _09963_/B vssd1 vssd1 vccd1 vccd1 _09963_/Y sky130_fd_sc_hd__nor2_1
X_05086_ _08956_/B vssd1 vssd1 vccd1 vccd1 _09538_/B sky130_fd_sc_hd__clkinv_2
XFILLER_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_65_wb_clk_i clkbuf_leaf_69_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11800_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08914_ _11316_/Q _08946_/B vssd1 vssd1 vccd1 vccd1 _08914_/X sky130_fd_sc_hd__or2_1
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _11715_/Q _09570_/A _09572_/D _11703_/Q _09893_/X vssd1 vssd1 vccd1 vccd1
+ _09899_/B sky130_fd_sc_hd__a221o_1
XFILLER_44_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _08847_/A _08845_/B vssd1 vssd1 vccd1 vccd1 _11280_/D sky130_fd_sc_hd__or2_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _11244_/Q _08804_/B vssd1 vssd1 vccd1 vccd1 _08776_/X sky130_fd_sc_hd__or2_1
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05988_ _05988_/A _05988_/B _05988_/C vssd1 vssd1 vccd1 vccd1 _05988_/X sky130_fd_sc_hd__and3_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07727_ _08789_/A1 _07755_/A2 _07726_/X _07205_/A vssd1 vssd1 vccd1 vccd1 _10664_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07658_ _10622_/Q _09214_/A _07663_/S vssd1 vssd1 vccd1 vccd1 _07659_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06609_ _10386_/Q _07939_/A _08286_/A _10727_/Q vssd1 vssd1 vccd1 vccd1 _06609_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07589_ _07076_/A _10578_/Q _07589_/S vssd1 vssd1 vccd1 vccd1 _07590_/B sky130_fd_sc_hd__mux2_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09328_ _11518_/Q _09326_/X _09327_/X vssd1 vssd1 vccd1 vccd1 _11518_/D sky130_fd_sc_hd__a21o_1
XFILLER_22_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09259_ _10168_/A1 _09249_/X _09258_/X _09267_/C1 vssd1 vssd1 vccd1 vccd1 _11482_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11221_ _11629_/CLK _11221_/D vssd1 vssd1 vccd1 vccd1 _11221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11152_ _11325_/CLK _11152_/D vssd1 vssd1 vccd1 vccd1 _11152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10103_ _10153_/A1 _10087_/X _10102_/X _10155_/C1 vssd1 vssd1 vccd1 vccd1 _11753_/D
+ sky130_fd_sc_hd__o211a_1
X_11083_ _11651_/CLK _11083_/D vssd1 vssd1 vccd1 vccd1 _11083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10034_ _11707_/Q _07104_/A _10051_/S vssd1 vssd1 vccd1 vccd1 _10035_/B sky130_fd_sc_hd__mux2_1
XFILLER_76_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10936_ _11023_/CLK _10936_/D vssd1 vssd1 vccd1 vccd1 _10936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10867_ _11485_/CLK _10867_/D vssd1 vssd1 vccd1 vccd1 _10867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _10798_/CLK _10798_/D vssd1 vssd1 vccd1 vccd1 _10798_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11419_ _11792_/CLK _11419_/D vssd1 vssd1 vccd1 vccd1 _11419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06960_ _09539_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09488_/C sky130_fd_sc_hd__nand2_4
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05911_ _10476_/Q _06803_/A2 _05910_/X _06997_/A vssd1 vssd1 vccd1 vccd1 _05911_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06891_ _06892_/A _06892_/B vssd1 vssd1 vccd1 vccd1 _07151_/C sky130_fd_sc_hd__nor2_8
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ _09237_/A0 _08621_/S _08629_/X _07003_/B vssd1 vssd1 vccd1 vccd1 _11169_/D
+ sky130_fd_sc_hd__o211a_1
X_05842_ _05833_/X _05834_/X _05836_/X _05841_/X vssd1 vssd1 vccd1 vccd1 _05842_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_95_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08561_ _11135_/Q _07048_/A _08577_/S vssd1 vssd1 vccd1 vccd1 _08562_/B sky130_fd_sc_hd__mux2_1
XFILLER_81_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05773_ _07690_/A _05767_/X _05772_/X _08243_/A _05762_/X vssd1 vssd1 vccd1 vccd1
+ _05773_/X sky130_fd_sc_hd__o311a_2
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07512_ _07916_/A _07512_/B vssd1 vssd1 vccd1 vccd1 _10540_/D sky130_fd_sc_hd__or2_1
XFILLER_23_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08492_ _08492_/A _08492_/B vssd1 vssd1 vccd1 vccd1 _11096_/D sky130_fd_sc_hd__or2_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_112_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11462_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07443_ _09193_/A _07535_/S vssd1 vssd1 vccd1 vccd1 _07443_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07374_ _07939_/A _08649_/B _07643_/C vssd1 vssd1 vccd1 vccd1 _07380_/S sky130_fd_sc_hd__and3_4
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09113_ _11403_/Q _09127_/B vssd1 vssd1 vccd1 vccd1 _09113_/X sky130_fd_sc_hd__or2_1
XFILLER_149_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06325_ _10826_/Q _07994_/A _06630_/B1 _11017_/Q _06324_/X vssd1 vssd1 vccd1 vccd1
+ _06325_/X sky130_fd_sc_hd__o221a_1
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ _11371_/Q _09038_/X _09043_/X vssd1 vssd1 vccd1 vccd1 _11371_/D sky130_fd_sc_hd__a21o_1
X_06256_ _11773_/Q _10119_/A vssd1 vssd1 vccd1 vccd1 _06256_/X sky130_fd_sc_hd__or2_1
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05207_ _10432_/Q _10431_/Q _05413_/S vssd1 vssd1 vccd1 vccd1 _05214_/B sky130_fd_sc_hd__mux2_2
XFILLER_89_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06187_ _11808_/Q _10180_/A _06185_/X _06186_/X vssd1 vssd1 vccd1 vccd1 _06187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05138_ _10636_/Q _10635_/Q _06939_/A vssd1 vssd1 vccd1 vccd1 _05140_/C sky130_fd_sc_hd__mux2_1
XFILLER_143_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout900 fanout901/X vssd1 vssd1 vccd1 vccd1 _06737_/A2 sky130_fd_sc_hd__buf_6
XFILLER_85_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout911 _07151_/A vssd1 vssd1 vccd1 vccd1 _07083_/B sky130_fd_sc_hd__buf_6
Xfanout922 _05092_/Y vssd1 vssd1 vccd1 vccd1 _06297_/C1 sky130_fd_sc_hd__buf_8
X_09946_ _10689_/Q _09573_/B _09573_/C _10373_/Q vssd1 vssd1 vccd1 vccd1 _09946_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout933 _10013_/A0 vssd1 vssd1 vccd1 vccd1 _10162_/A1 sky130_fd_sc_hd__buf_6
Xfanout944 _08647_/A vssd1 vssd1 vccd1 vccd1 _10135_/A0 sky130_fd_sc_hd__buf_6
Xfanout955 _09234_/A0 vssd1 vssd1 vccd1 vccd1 _09182_/A0 sky130_fd_sc_hd__buf_6
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout966 _08933_/A1 vssd1 vssd1 vccd1 vccd1 _08846_/A0 sky130_fd_sc_hd__buf_8
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout977 _10181_/A0 vssd1 vssd1 vccd1 vccd1 _10088_/A1 sky130_fd_sc_hd__buf_6
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _10561_/Q _09877_/A2 _09877_/B1 _10562_/Q _09876_/X vssd1 vssd1 vccd1 vccd1
+ _09880_/C sky130_fd_sc_hd__a221o_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout988 _11870_/A vssd1 vssd1 vccd1 vccd1 _07297_/A sky130_fd_sc_hd__buf_6
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout999 _06357_/C1 vssd1 vssd1 vccd1 vccd1 _06670_/D1 sky130_fd_sc_hd__buf_12
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08828_ _11272_/Q _08840_/B vssd1 vssd1 vccd1 vccd1 _08828_/X sky130_fd_sc_hd__or2_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _08661_/A _08760_/S _08758_/X _09267_/C1 vssd1 vssd1 vccd1 vccd1 _11236_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11770_ _11770_/CLK _11770_/D vssd1 vssd1 vccd1 vccd1 _11770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10798_/CLK _10721_/D vssd1 vssd1 vccd1 vccd1 _10721_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10652_ _11151_/CLK _10652_/D vssd1 vssd1 vccd1 vccd1 _10652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10583_ _11628_/CLK _10583_/D vssd1 vssd1 vccd1 vccd1 _10583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11204_ _11329_/CLK _11204_/D vssd1 vssd1 vccd1 vccd1 _11204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11135_ _11224_/CLK _11135_/D vssd1 vssd1 vccd1 vccd1 _11135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11066_ _11067_/CLK _11066_/D vssd1 vssd1 vccd1 vccd1 _11066_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10017_ _10017_/A0 _11699_/Q _10028_/B vssd1 vssd1 vccd1 vccd1 _10018_/B sky130_fd_sc_hd__mux2_1
XFILLER_92_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10919_ _11770_/CLK _10919_/D vssd1 vssd1 vccd1 vccd1 _10919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06110_ _10559_/Q _07540_/A _06805_/B1 _10535_/Q vssd1 vssd1 vccd1 vccd1 _06110_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_69_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07090_ _07090_/A _07318_/A vssd1 vssd1 vccd1 vccd1 _07090_/X sky130_fd_sc_hd__or2_4
XFILLER_133_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06041_ _10685_/Q _06370_/A2 _07819_/A _10719_/Q vssd1 vssd1 vccd1 vccd1 _06041_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_114_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09800_ _10525_/Q _09565_/B _09948_/B1 _10290_/Q _09799_/X vssd1 vssd1 vccd1 vccd1
+ _09815_/A sky130_fd_sc_hd__a221o_1
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout218 _07353_/Y vssd1 vssd1 vccd1 vccd1 _07355_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_113_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout229 _07188_/S vssd1 vssd1 vccd1 vccd1 _07123_/B1 sky130_fd_sc_hd__clkbuf_2
X_07992_ _08578_/A _07992_/B vssd1 vssd1 vccd1 vccd1 _10821_/D sky130_fd_sc_hd__and2_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09731_ _09731_/A _09731_/B _09731_/C _09731_/D vssd1 vssd1 vccd1 vccd1 _09739_/A
+ sky130_fd_sc_hd__or4_1
X_06943_ _05473_/B _09553_/A vssd1 vssd1 vccd1 vccd1 _06944_/A sky130_fd_sc_hd__and2b_2
XFILLER_101_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09662_ _11630_/Q _09660_/Y _09661_/X _09641_/Y _09959_/A vssd1 vssd1 vccd1 vccd1
+ _11630_/D sky130_fd_sc_hd__a221o_1
XFILLER_67_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06874_ _10769_/Q _07854_/A vssd1 vssd1 vccd1 vccd1 _06874_/X sky130_fd_sc_hd__or2_1
XFILLER_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08613_ _09101_/A1 _11161_/Q _08623_/S vssd1 vssd1 vccd1 vccd1 _08614_/B sky130_fd_sc_hd__mux2_1
X_05825_ _11747_/Q _05953_/A2 _06214_/B1 _11783_/Q _06349_/C1 vssd1 vssd1 vccd1 vccd1
+ _05825_/X sky130_fd_sc_hd__o221a_1
X_09593_ _09593_/A _09593_/B _09593_/C _09593_/D vssd1 vssd1 vccd1 vccd1 _09594_/D
+ sky130_fd_sc_hd__nor4_2
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08544_ _08893_/A1 _08506_/X _08543_/X _08919_/C1 vssd1 vssd1 vccd1 vccd1 _11121_/D
+ sky130_fd_sc_hd__o211a_1
X_05756_ _11676_/Q _08594_/A _05752_/X _05755_/X vssd1 vssd1 vccd1 vccd1 _05762_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08475_ _11088_/Q _08503_/B vssd1 vssd1 vccd1 vccd1 _08475_/X sky130_fd_sc_hd__or2_1
XFILLER_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05687_ _11162_/Q _05524_/Y _05585_/Y _11166_/Q vssd1 vssd1 vccd1 vccd1 _05687_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07426_ _10026_/A _07426_/B vssd1 vssd1 vccd1 vccd1 _10489_/D sky130_fd_sc_hd__or2_1
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07357_ _07235_/X _10450_/Q _07357_/S vssd1 vssd1 vccd1 vccd1 _10450_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06308_ _10286_/Q _06308_/A2 _06373_/B1 _10317_/Q _06305_/X vssd1 vssd1 vccd1 vccd1
+ _06309_/C sky130_fd_sc_hd__o221a_2
X_07288_ _10051_/A1 _09187_/S _07287_/X _07902_/C1 vssd1 vssd1 vccd1 vccd1 _10412_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_wb_clk_i clkbuf_leaf_85_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11572_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_152_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09027_ _11364_/Q _09035_/B vssd1 vssd1 vccd1 vccd1 _09027_/X sky130_fd_sc_hd__or2_1
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06239_ _10285_/Q _06308_/A2 _06235_/X _06238_/X vssd1 vssd1 vccd1 vccd1 _06239_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_151_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout730 _06728_/B1 vssd1 vssd1 vccd1 vccd1 _06805_/B1 sky130_fd_sc_hd__buf_6
Xfanout741 _05750_/Y vssd1 vssd1 vccd1 vccd1 _09292_/A sky130_fd_sc_hd__buf_12
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout752 _08994_/A vssd1 vssd1 vccd1 vccd1 _10137_/A sky130_fd_sc_hd__buf_4
X_09929_ input7/X _09889_/Y _09926_/Y vssd1 vssd1 vccd1 vccd1 _09929_/X sky130_fd_sc_hd__a21o_1
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout763 _06739_/A2 vssd1 vssd1 vccd1 vccd1 _06718_/B1 sky130_fd_sc_hd__buf_4
XFILLER_63_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout774 _08300_/A vssd1 vssd1 vccd1 vccd1 _06628_/B1 sky130_fd_sc_hd__buf_6
Xfanout785 _06806_/A2 vssd1 vssd1 vccd1 vccd1 _06877_/B1 sky130_fd_sc_hd__buf_6
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout796 _06152_/B vssd1 vssd1 vccd1 vccd1 _06636_/A2 sky130_fd_sc_hd__buf_6
XFILLER_59_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _09571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _09976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _07104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _10017_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _05737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_156 _07105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_167 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11753_ _11791_/CLK _11753_/D vssd1 vssd1 vccd1 vccd1 _11753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_178 _06674_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_189 _07059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10765_/CLK _10704_/D vssd1 vssd1 vccd1 vccd1 _10704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11684_ _11684_/CLK _11684_/D vssd1 vssd1 vccd1 vccd1 _11684_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10635_ _10644_/CLK _10635_/D vssd1 vssd1 vccd1 vccd1 _10635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10566_ _11472_/CLK _10566_/D vssd1 vssd1 vccd1 vccd1 _10566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10497_ _10804_/CLK _10497_/D vssd1 vssd1 vccd1 vccd1 _10497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11118_ _11329_/CLK _11118_/D vssd1 vssd1 vccd1 vccd1 _11118_/Q sky130_fd_sc_hd__dfxtp_1
X_11049_ _11575_/CLK _11049_/D vssd1 vssd1 vccd1 vccd1 _11049_/Q sky130_fd_sc_hd__dfxtp_1
Xinput7 ram_val_in[1] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_4
XFILLER_64_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05610_ _09552_/A1 _11397_/Q _11391_/Q _05078_/A vssd1 vssd1 vccd1 vccd1 _05610_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06590_ _06586_/X _06589_/X _07689_/A _06584_/X vssd1 vssd1 vccd1 vccd1 _06590_/X
+ sky130_fd_sc_hd__a211o_2
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05541_ _05631_/A2 _11358_/Q _11354_/Q _05631_/B1 _05539_/X vssd1 vssd1 vccd1 vccd1
+ _05541_/X sky130_fd_sc_hd__a221o_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08260_ _10962_/Q _08284_/B vssd1 vssd1 vccd1 vccd1 _08260_/X sky130_fd_sc_hd__or2_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05472_ _09681_/A _05472_/B vssd1 vssd1 vccd1 vccd1 _05473_/B sky130_fd_sc_hd__or2_2
X_07211_ _07211_/A _07420_/A vssd1 vssd1 vccd1 vccd1 _07211_/X sky130_fd_sc_hd__or2_1
X_08191_ _10930_/Q _08197_/S _07644_/Y _07098_/B vssd1 vssd1 vccd1 vccd1 _10930_/D
+ sky130_fd_sc_hd__o22a_1
X_07142_ _10332_/Q _07145_/B _07188_/S _07141_/X vssd1 vssd1 vccd1 vccd1 _10332_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07073_ _10047_/A1 _07074_/S _07072_/X _07147_/B vssd1 vssd1 vccd1 vccd1 _10295_/D
+ sky130_fd_sc_hd__o211a_1
X_06024_ _11383_/Q _08383_/A _06219_/A2 _11393_/Q _06023_/X vssd1 vssd1 vccd1 vccd1
+ _06024_/X sky130_fd_sc_hd__o221a_1
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07975_ _10811_/Q _07010_/A _07991_/S vssd1 vssd1 vccd1 vccd1 _07976_/B sky130_fd_sc_hd__mux2_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06926_ _10110_/A0 _10204_/Q _06934_/S vssd1 vssd1 vccd1 vccd1 _10204_/D sky130_fd_sc_hd__mux2_1
X_09714_ _10412_/Q _09882_/B1 _09567_/D _10406_/Q vssd1 vssd1 vccd1 vccd1 _09714_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06857_ _10362_/Q _06872_/A2 _06857_/B1 _11722_/Q vssd1 vssd1 vccd1 vccd1 _06857_/X
+ sky130_fd_sc_hd__o22a_1
X_09645_ _10310_/Q _09566_/A _09568_/C _10322_/Q _09644_/X vssd1 vssd1 vccd1 vccd1
+ _09650_/B sky130_fd_sc_hd__a221o_1
XFILLER_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05808_ _10869_/Q _07994_/A _06453_/B1 _10985_/Q vssd1 vssd1 vccd1 vccd1 _05808_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _09576_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09594_/B sky130_fd_sc_hd__or2_1
XFILLER_110_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ _10734_/Q _06710_/B _06787_/X _06849_/C1 vssd1 vssd1 vccd1 vccd1 _06788_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08527_ _08876_/A0 _11113_/Q _08529_/S vssd1 vssd1 vccd1 vccd1 _08528_/B sky130_fd_sc_hd__mux2_1
X_05739_ _05749_/A _11868_/A _05745_/A vssd1 vssd1 vccd1 vccd1 _05739_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_54_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08458_ _11079_/Q _08459_/S _07628_/S _07333_/B vssd1 vssd1 vccd1 vccd1 _11079_/D
+ sky130_fd_sc_hd__o22a_1
X_07409_ _07018_/A _10481_/Q _07425_/S vssd1 vssd1 vccd1 vccd1 _07410_/B sky130_fd_sc_hd__mux2_1
XFILLER_156_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08389_ _09364_/A1 _08414_/S _08388_/X _09168_/C1 vssd1 vssd1 vccd1 vccd1 _11035_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10420_ _10644_/CLK _10420_/D vssd1 vssd1 vccd1 vccd1 _10420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10351_ _10548_/CLK _10351_/D vssd1 vssd1 vccd1 vccd1 _10351_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10282_ _11766_/CLK _10282_/D vssd1 vssd1 vccd1 vccd1 _10282_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_105_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout560 fanout565/X vssd1 vssd1 vccd1 vccd1 _08618_/A sky130_fd_sc_hd__buf_4
XFILLER_120_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout571 _08781_/A vssd1 vssd1 vccd1 vccd1 _08682_/A sky130_fd_sc_hd__buf_2
Xfanout582 _05818_/Y vssd1 vssd1 vccd1 vccd1 _08970_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout593 _09403_/Y vssd1 vssd1 vccd1 vccd1 _09554_/B sky130_fd_sc_hd__buf_6
XFILLER_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _11809_/CLK _11805_/D vssd1 vssd1 vccd1 vccd1 _11805_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11736_ _11765_/CLK _11736_/D vssd1 vssd1 vccd1 vccd1 _11736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ _11735_/CLK _11667_/D vssd1 vssd1 vccd1 vccd1 _11667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10618_ _11310_/CLK _10618_/D vssd1 vssd1 vccd1 vccd1 _10618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11598_ _11650_/CLK _11598_/D vssd1 vssd1 vccd1 vccd1 _11598_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10549_ _10769_/CLK _10549_/D vssd1 vssd1 vccd1 vccd1 _10549_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_155_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07760_ _10681_/Q _07760_/B vssd1 vssd1 vccd1 vccd1 _07760_/X sky130_fd_sc_hd__or2_1
XFILLER_110_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06711_ _10390_/Q _06871_/A2 _06856_/A2 _10327_/Q _06710_/X vssd1 vssd1 vccd1 vccd1
+ _06711_/X sky130_fd_sc_hd__o221a_1
X_07691_ _08649_/A _08649_/C _09037_/C vssd1 vssd1 vccd1 vccd1 _08591_/B sky130_fd_sc_hd__and3_4
XFILLER_38_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09430_ _11631_/Q _09430_/B vssd1 vssd1 vccd1 vccd1 _09672_/B sky130_fd_sc_hd__nand2_8
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06642_ _10473_/Q _06642_/A2 _06641_/X _06642_/C1 vssd1 vssd1 vccd1 vccd1 _06642_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09361_ _10161_/A1 _09359_/X _09360_/X _09995_/C1 vssd1 vssd1 vccd1 vccd1 _11538_/D
+ sky130_fd_sc_hd__o211a_1
X_06573_ _11116_/Q _06646_/A2 _06571_/X _06572_/X vssd1 vssd1 vccd1 vccd1 _06573_/X
+ sky130_fd_sc_hd__a211o_1
X_08312_ _09999_/A0 _10991_/Q _08321_/S vssd1 vssd1 vccd1 vccd1 _10991_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11233_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05524_ _05524_/A _05524_/B vssd1 vssd1 vccd1 vccd1 _05524_/Y sky130_fd_sc_hd__nor2_8
XFILLER_21_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09292_ _09292_/A _10158_/B _10158_/C vssd1 vssd1 vccd1 vccd1 _09310_/B sky130_fd_sc_hd__and3_4
XFILLER_21_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _05737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_23 _06761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _08243_/A _08243_/B _08243_/C _08243_/D vssd1 vssd1 vccd1 vccd1 _08243_/X
+ sky130_fd_sc_hd__or4_4
XANTENNA_34 _08545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05455_ _10769_/Q _09953_/B1 _09884_/A2 _10807_/Q _05454_/X vssd1 vssd1 vccd1 vccd1
+ _05469_/A sky130_fd_sc_hd__a221o_1
XFILLER_53_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_45 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_56 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 _11615_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ _07018_/A _10916_/Q _08182_/S vssd1 vssd1 vccd1 vccd1 _10916_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05386_ _10471_/Q _10470_/Q _05397_/S vssd1 vssd1 vccd1 vccd1 _05389_/B sky130_fd_sc_hd__mux2_1
XANTENNA_89 _08441_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07125_ _10322_/Q _07126_/B _07186_/S _08817_/B2 vssd1 vssd1 vccd1 vccd1 _10322_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07056_ _10286_/Q _07047_/B _07490_/S _07022_/B vssd1 vssd1 vccd1 vccd1 _10286_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput130 _11610_/Q vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_4
Xoutput141 _11621_/Q vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__buf_4
XFILLER_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput152 _11575_/Q vssd1 vssd1 vccd1 vccd1 ram_addr[6] sky130_fd_sc_hd__buf_4
X_06007_ _11026_/Q _06629_/A2 _06453_/B1 _10636_/Q vssd1 vssd1 vccd1 vccd1 _06007_/X
+ sky130_fd_sc_hd__o22a_1
Xoutput163 _11583_/Q vssd1 vssd1 vccd1 vccd1 rom_addr[5] sky130_fd_sc_hd__buf_4
XFILLER_115_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput174 _11872_/X vssd1 vssd1 vccd1 vccd1 wb_rom_adrb[6] sky130_fd_sc_hd__buf_4
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput185 _05491_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_4
Xoutput196 _05501_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_4
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07958_ _07070_/A _07820_/B _07821_/A _10800_/Q _07333_/A vssd1 vssd1 vccd1 vccd1
+ _10800_/D sky130_fd_sc_hd__a221o_1
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06909_ _10111_/A0 _06903_/X _06908_/X _06996_/C1 vssd1 vssd1 vccd1 vccd1 _10195_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07889_ _10763_/Q _07901_/B vssd1 vssd1 vccd1 vccd1 _07889_/X sky130_fd_sc_hd__or2_1
XFILLER_29_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09628_ _10718_/Q _09566_/B _09573_/B _10723_/Q vssd1 vssd1 vccd1 vccd1 _09628_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09559_ _11660_/Q _11645_/Q vssd1 vssd1 vccd1 vccd1 _09600_/B sky130_fd_sc_hd__and2_2
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ _11683_/CLK _11521_/D vssd1 vssd1 vccd1 vccd1 _11521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11452_ _11471_/CLK _11452_/D vssd1 vssd1 vccd1 vccd1 _11452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10403_ _10808_/CLK _10403_/D vssd1 vssd1 vccd1 vccd1 _10403_/Q sky130_fd_sc_hd__dfxtp_1
X_11383_ _11428_/CLK _11383_/D vssd1 vssd1 vccd1 vccd1 _11383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10334_ _11720_/CLK _10334_/D vssd1 vssd1 vccd1 vccd1 _10334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _11810_/CLK _10265_/D vssd1 vssd1 vccd1 vccd1 _10265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10196_ _11755_/CLK _10196_/D vssd1 vssd1 vccd1 vccd1 _10196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout390 _07599_/A vssd1 vssd1 vccd1 vccd1 _07617_/A sky130_fd_sc_hd__buf_6
XFILLER_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11719_ _11719_/CLK _11719_/D vssd1 vssd1 vccd1 vccd1 _11719_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05240_ _05085_/Y _10864_/Q _10787_/Q _09444_/A _05239_/X vssd1 vssd1 vccd1 vccd1
+ _05248_/A sky130_fd_sc_hd__a221o_2
XFILLER_147_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 rom_value[0] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_2
XFILLER_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput21 rom_value[1] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
Xinput32 rom_value[2] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_2
Xinput43 wb_rom_val[10] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_2
XFILLER_128_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput54 wb_rom_val[20] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_4
X_05171_ _11230_/Q _11229_/Q _05349_/S vssd1 vssd1 vccd1 vccd1 _05178_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput65 wb_rom_val[30] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_4
Xinput76 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_4
Xinput87 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_137_wb_clk_i clkbuf_4_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10255_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput98 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08930_ _11324_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08930_/X sky130_fd_sc_hd__or2_1
XFILLER_130_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08861_ _08873_/A _08861_/B vssd1 vssd1 vccd1 vccd1 _11287_/D sky130_fd_sc_hd__or2_1
XFILLER_44_1338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07812_ _07812_/A _07812_/B vssd1 vssd1 vccd1 vccd1 _10713_/D sky130_fd_sc_hd__or2_1
X_08792_ _08883_/A1 _11252_/Q _08792_/S vssd1 vssd1 vccd1 vccd1 _08793_/B sky130_fd_sc_hd__mux2_1
XFILLER_85_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07743_ _08423_/A1 _07761_/A2 _07742_/X _07932_/C1 vssd1 vssd1 vccd1 vccd1 _10672_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07674_ _08655_/B _08663_/S vssd1 vssd1 vccd1 vccd1 _07674_/X sky130_fd_sc_hd__or2_4
XFILLER_65_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _11334_/Q _11574_/Q _09414_/S vssd1 vssd1 vccd1 vccd1 _11574_/D sky130_fd_sc_hd__mux2_1
X_06625_ _10868_/Q _06976_/A _06903_/A _10908_/Q vssd1 vssd1 vccd1 vccd1 _06625_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_34_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09344_ _09995_/A1 _09326_/X _09343_/X _09993_/C1 vssd1 vssd1 vccd1 vccd1 _11526_/D
+ sky130_fd_sc_hd__o211a_1
X_06556_ _10850_/Q _06643_/A2 _06556_/B1 _11084_/Q _06555_/X vssd1 vssd1 vccd1 vccd1
+ _06556_/X sky130_fd_sc_hd__o221a_1
XFILLER_40_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05507_ _10252_/Q input65/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05507_/X sky130_fd_sc_hd__mux2_4
XFILLER_51_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09275_ _09275_/A1 _09271_/X _09274_/X _09289_/C1 vssd1 vssd1 vccd1 vccd1 _11489_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06487_ _11324_/Q _06648_/A2 _09131_/A _11296_/Q _08243_/B vssd1 vssd1 vccd1 vccd1
+ _06487_/X sky130_fd_sc_hd__a221o_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08226_ _08839_/A _08226_/B vssd1 vssd1 vccd1 vccd1 _10947_/D sky130_fd_sc_hd__or2_1
X_05438_ _10664_/Q _09947_/A2 _09568_/B _10657_/Q vssd1 vssd1 vccd1 vccd1 _05438_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_101_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08157_ _10172_/A1 _08162_/S _08156_/X _07011_/B vssd1 vssd1 vccd1 vccd1 _10904_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05369_ _10829_/Q _10828_/Q _05430_/S vssd1 vssd1 vccd1 vccd1 _05373_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07108_ _07333_/A _07335_/B vssd1 vssd1 vccd1 vccd1 _07108_/X sky130_fd_sc_hd__or2_4
XFILLER_107_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08088_ _07303_/X _08015_/S _08087_/X _08427_/A vssd1 vssd1 vccd1 vccd1 _10869_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07039_ _07039_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _07040_/B sky130_fd_sc_hd__and2_4
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10050_ _10050_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _11716_/D sky130_fd_sc_hd__or2_1
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10952_ _11234_/CLK _10952_/D vssd1 vssd1 vccd1 vccd1 _10952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10883_ _11776_/CLK _10883_/D vssd1 vssd1 vccd1 vccd1 _10883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11504_ _11800_/CLK _11504_/D vssd1 vssd1 vccd1 vccd1 _11504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ _11473_/CLK _11435_/D vssd1 vssd1 vccd1 vccd1 _11435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11366_ _11366_/CLK _11366_/D vssd1 vssd1 vccd1 vccd1 _11366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10317_ _10812_/CLK _10317_/D vssd1 vssd1 vccd1 vccd1 _10317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ _11325_/CLK _11297_/D vssd1 vssd1 vccd1 vccd1 _11297_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10248_ _11712_/CLK _10248_/D vssd1 vssd1 vccd1 vccd1 _10248_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10179_ _11801_/Q _10159_/X _10178_/X vssd1 vssd1 vccd1 vccd1 _11801_/D sky130_fd_sc_hd__a21o_1
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06410_ _10425_/Q _06541_/A2 _06538_/B1 _10643_/Q vssd1 vssd1 vccd1 vccd1 _06410_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07390_ _10471_/Q _07393_/S _07655_/S _08817_/B2 vssd1 vssd1 vccd1 vccd1 _10471_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06341_ _06535_/A _06317_/X _06339_/X _06340_/X vssd1 vssd1 vccd1 vccd1 _06341_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_148_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09060_ _09060_/A _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09060_/X sky130_fd_sc_hd__or3_4
X_06272_ _07151_/B _06245_/X _06250_/X _06234_/X vssd1 vssd1 vccd1 vccd1 _06272_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_148_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08011_ _10132_/A0 _10830_/Q _08011_/S vssd1 vssd1 vccd1 vccd1 _08012_/B sky130_fd_sc_hd__mux2_1
X_05223_ _05223_/A _05223_/B _05223_/C _05223_/D vssd1 vssd1 vccd1 vccd1 _05224_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_116_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05154_ _10948_/Q _10947_/Q _09680_/B vssd1 vssd1 vccd1 vccd1 _05156_/C sky130_fd_sc_hd__mux2_1
X_09962_ _11664_/Q _09823_/Y _09963_/B vssd1 vssd1 vccd1 vccd1 _11664_/D sky130_fd_sc_hd__mux2_1
X_05085_ _05326_/S vssd1 vssd1 vccd1 vccd1 _05085_/Y sky130_fd_sc_hd__inv_4
XFILLER_143_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08913_ _09276_/A1 _08945_/A2 _08912_/X _09078_/C1 vssd1 vssd1 vccd1 vccd1 _11315_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09893_ _11745_/Q _09572_/A _09571_/C _11717_/Q vssd1 vssd1 vccd1 vccd1 _09893_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08844_ _10171_/A1 _11280_/Q _08850_/S vssd1 vssd1 vccd1 vccd1 _08845_/B sky130_fd_sc_hd__mux2_1
XFILLER_111_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08775_ _08793_/A _08775_/B vssd1 vssd1 vccd1 vccd1 _11243_/D sky130_fd_sc_hd__or2_1
X_05987_ _11106_/Q _06737_/A2 _08765_/A _11242_/Q vssd1 vssd1 vccd1 vccd1 _05988_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11733_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07726_ _10664_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07726_/X sky130_fd_sc_hd__or2_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07657_ _10621_/Q _07663_/S _07246_/S _07052_/X vssd1 vssd1 vccd1 vccd1 _10621_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06608_ _10368_/Q _09358_/A _09976_/A _10272_/Q _07151_/A vssd1 vssd1 vccd1 vccd1
+ _06608_/X sky130_fd_sc_hd__a221o_1
X_07588_ _07926_/A _07588_/B vssd1 vssd1 vccd1 vccd1 _10577_/D sky130_fd_sc_hd__or2_1
XFILLER_129_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09327_ _10161_/A1 _09343_/B _08618_/A vssd1 vssd1 vccd1 vccd1 _09327_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06539_ _11282_/Q _06539_/A2 _06539_/B1 _10596_/Q _06624_/C1 vssd1 vssd1 vccd1 vccd1
+ _06539_/X sky130_fd_sc_hd__o221a_2
XFILLER_107_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ _11482_/Q _09266_/B vssd1 vssd1 vccd1 vccd1 _09258_/X sky130_fd_sc_hd__or2_1
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08209_ _10939_/Q _08902_/C vssd1 vssd1 vccd1 vccd1 _08209_/X sky130_fd_sc_hd__or2_1
X_09189_ _11440_/Q _09175_/Y _09176_/Y _07043_/X vssd1 vssd1 vccd1 vccd1 _11440_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11220_ _11220_/CLK _11220_/D vssd1 vssd1 vccd1 vccd1 _11220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11151_ _11151_/CLK _11151_/D vssd1 vssd1 vccd1 vccd1 _11151_/Q sky130_fd_sc_hd__dfxtp_1
X_10102_ _11753_/Q _10104_/B vssd1 vssd1 vccd1 vccd1 _10102_/X sky130_fd_sc_hd__or2_1
XFILLER_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11082_ _11140_/CLK _11082_/D vssd1 vssd1 vccd1 vccd1 _11082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10033_ _10039_/A _10033_/B vssd1 vssd1 vccd1 vccd1 _11706_/D sky130_fd_sc_hd__or2_1
XFILLER_153_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10935_ _11023_/CLK _10935_/D vssd1 vssd1 vccd1 vccd1 _10935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10866_ _11235_/CLK _10866_/D vssd1 vssd1 vccd1 vccd1 _10866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10797_ _10981_/CLK _10797_/D vssd1 vssd1 vccd1 vccd1 _10797_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11418_ _11792_/CLK _11418_/D vssd1 vssd1 vccd1 vccd1 _11418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11349_ _11485_/CLK _11349_/D vssd1 vssd1 vccd1 vccd1 _11349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05910_ _10683_/Q _07904_/A _07539_/A _10312_/Q _05909_/X vssd1 vssd1 vccd1 vccd1
+ _05910_/X sky130_fd_sc_hd__o221a_1
X_06890_ input76/X _10255_/D vssd1 vssd1 vccd1 vccd1 _06890_/Y sky130_fd_sc_hd__nand2_4
X_05841_ _10204_/Q _10072_/A _05837_/X _05840_/X vssd1 vssd1 vccd1 vccd1 _05841_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05772_ _10203_/Q _06351_/A2 _05768_/X _05771_/X vssd1 vssd1 vccd1 vccd1 _05772_/X
+ sky130_fd_sc_hd__o211a_1
X_08560_ _08560_/A _08649_/B _08560_/C vssd1 vssd1 vccd1 vccd1 _08567_/S sky130_fd_sc_hd__and3_2
XFILLER_78_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07511_ _08931_/A1 _10540_/Q _07513_/S vssd1 vssd1 vccd1 vccd1 _07512_/B sky130_fd_sc_hd__mux2_1
X_08491_ _10118_/A0 _11096_/Q _08497_/S vssd1 vssd1 vccd1 vccd1 _08492_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07442_ _09227_/A _07513_/S vssd1 vssd1 vccd1 vccd1 _07442_/Y sky130_fd_sc_hd__nand2_2
XFILLER_62_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07373_ _10461_/Q _08901_/A1 _07373_/S vssd1 vssd1 vccd1 vccd1 _10461_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09112_ _11402_/Q _09110_/X _09111_/X vssd1 vssd1 vccd1 vccd1 _11402_/D sky130_fd_sc_hd__a21o_1
X_06324_ _10650_/Q _07692_/A _06632_/A2 _10893_/Q vssd1 vssd1 vccd1 vccd1 _06324_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_149_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09043_ _09276_/A1 _09055_/B _09173_/B1 vssd1 vssd1 vccd1 vccd1 _09043_/X sky130_fd_sc_hd__a21o_1
XFILLER_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06255_ _06255_/A _06255_/B _06255_/C vssd1 vssd1 vccd1 vccd1 _06255_/X sky130_fd_sc_hd__and3_1
X_05206_ _09444_/A _10901_/Q _10430_/Q _05085_/Y _05205_/X vssd1 vssd1 vccd1 vccd1
+ _05214_/A sky130_fd_sc_hd__a221o_2
XFILLER_135_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06186_ _10262_/Q _06976_/A _06903_/A _10199_/Q vssd1 vssd1 vccd1 vccd1 _06186_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_102_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05137_ _10640_/Q _10639_/Q _05414_/S vssd1 vssd1 vccd1 vccd1 _05140_/B sky130_fd_sc_hd__mux2_1
XFILLER_137_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout901 _05739_/Y vssd1 vssd1 vccd1 vccd1 fanout901/X sky130_fd_sc_hd__buf_8
XFILLER_137_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout912 _07151_/A vssd1 vssd1 vccd1 vccd1 _06642_/C1 sky130_fd_sc_hd__buf_4
X_09945_ _10688_/Q _09571_/B _09572_/D _10365_/Q vssd1 vssd1 vccd1 vccd1 _09945_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout923 _06189_/A1 vssd1 vssd1 vccd1 vccd1 _07083_/A sky130_fd_sc_hd__buf_8
Xfanout934 input99/X vssd1 vssd1 vccd1 vccd1 _10013_/A0 sky130_fd_sc_hd__buf_6
Xfanout945 input94/X vssd1 vssd1 vccd1 vccd1 _08647_/A sky130_fd_sc_hd__buf_4
XFILLER_86_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout956 _09234_/A0 vssd1 vssd1 vccd1 vccd1 _08937_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout967 input91/X vssd1 vssd1 vccd1 vccd1 _08933_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09876_ _10578_/Q _09876_/A2 _09876_/B1 _10564_/Q vssd1 vssd1 vccd1 vccd1 _09876_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout978 _08669_/A0 vssd1 vssd1 vccd1 vccd1 _10181_/A0 sky130_fd_sc_hd__buf_8
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout989 input83/X vssd1 vssd1 vccd1 vccd1 _11870_/A sky130_fd_sc_hd__buf_12
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08839_/A _08827_/B vssd1 vssd1 vccd1 vccd1 _11271_/D sky130_fd_sc_hd__or2_1
XFILLER_73_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _11236_/Q _08762_/B vssd1 vssd1 vccd1 vccd1 _08758_/X sky130_fd_sc_hd__or2_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _10013_/A0 _07755_/A2 _07708_/X _07868_/C1 vssd1 vssd1 vccd1 vccd1 _10655_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _08876_/A0 _11199_/Q _08707_/S vssd1 vssd1 vccd1 vccd1 _08690_/B sky130_fd_sc_hd__mux2_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10720_ _11713_/CLK _10720_/D vssd1 vssd1 vccd1 vccd1 _10720_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10651_ _11270_/CLK _10651_/D vssd1 vssd1 vccd1 vccd1 _10651_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10582_ _11280_/CLK _10582_/D vssd1 vssd1 vccd1 vccd1 _10582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11203_ _11329_/CLK _11203_/D vssd1 vssd1 vccd1 vccd1 _11203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11134_ _11268_/CLK _11134_/D vssd1 vssd1 vccd1 vccd1 _11134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11065_ _11067_/CLK _11065_/D vssd1 vssd1 vccd1 vccd1 _11065_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10016_ _10026_/A _10016_/B vssd1 vssd1 vccd1 vccd1 _11698_/D sky130_fd_sc_hd__or2_1
XFILLER_37_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10918_ _11779_/CLK _10918_/D vssd1 vssd1 vccd1 vccd1 _10918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10849_ _11140_/CLK _10849_/D vssd1 vssd1 vccd1 vccd1 _10849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06040_ _10382_/Q _06871_/A2 _06999_/A _10508_/Q vssd1 vssd1 vccd1 vccd1 _06040_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout219 _07353_/Y vssd1 vssd1 vccd1 vccd1 _07357_/S sky130_fd_sc_hd__buf_2
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07991_ _10821_/Q _10135_/A0 _07991_/S vssd1 vssd1 vccd1 vccd1 _07992_/B sky130_fd_sc_hd__mux2_1
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09730_ _11472_/Q _09876_/A2 _09573_/A _11467_/Q _09729_/X vssd1 vssd1 vccd1 vccd1
+ _09731_/D sky130_fd_sc_hd__a221o_1
X_06942_ _06942_/A _06942_/B _11599_/Q _06945_/B vssd1 vssd1 vccd1 vccd1 _09668_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09661_ _09660_/Y _09661_/B vssd1 vssd1 vccd1 vccd1 _09661_/X sky130_fd_sc_hd__and2b_1
XFILLER_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06873_ _10532_/Q _06873_/A2 _06870_/X _06872_/X _06873_/D1 vssd1 vssd1 vccd1 vccd1
+ _06873_/X sky130_fd_sc_hd__o2111a_1
XFILLER_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08612_ _08847_/A _08612_/B vssd1 vssd1 vccd1 vccd1 _11160_/D sky130_fd_sc_hd__or2_1
X_05824_ _11519_/Q _09326_/A _06363_/A2 _11479_/Q _05823_/X vssd1 vssd1 vccd1 vccd1
+ _05824_/X sky130_fd_sc_hd__o221a_1
X_09592_ _10512_/Q _09947_/A2 _09573_/B _10511_/Q _09579_/X vssd1 vssd1 vccd1 vccd1
+ _09593_/D sky130_fd_sc_hd__a221o_1
XFILLER_55_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05755_ _11538_/Q _09359_/A _05753_/X _05754_/X vssd1 vssd1 vccd1 vccd1 _05755_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08543_ _11121_/Q _08545_/B vssd1 vssd1 vccd1 vccd1 _08543_/X sky130_fd_sc_hd__or2_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05686_ _11163_/Q _05555_/Y _05627_/Y _11152_/Q _05685_/X vssd1 vssd1 vccd1 vccd1
+ _05691_/A sky130_fd_sc_hd__a221o_1
X_08474_ _10088_/A1 _08497_/S _08473_/X _09022_/C1 vssd1 vssd1 vccd1 vccd1 _11087_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07425_ _07031_/A _10489_/Q _07425_/S vssd1 vssd1 vccd1 vccd1 _07426_/B sky130_fd_sc_hd__mux2_1
XFILLER_126_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07356_ _07108_/X _10449_/Q _07357_/S vssd1 vssd1 vccd1 vccd1 _10449_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06307_ _10482_/Q _06803_/A2 _06857_/B1 _11703_/Q _06997_/A vssd1 vssd1 vccd1 vccd1
+ _06309_/B sky130_fd_sc_hd__o221a_1
X_07287_ _10412_/Q _09175_/B vssd1 vssd1 vccd1 vccd1 _07287_/X sky130_fd_sc_hd__or2_1
X_09026_ _10185_/A0 _09016_/X _09025_/X _09032_/C1 vssd1 vssd1 vccd1 vccd1 _11363_/D
+ sky130_fd_sc_hd__o211a_1
X_06238_ _10481_/Q _06238_/A2 _06237_/X _11869_/A vssd1 vssd1 vccd1 vccd1 _06238_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06169_ _11752_/Q _06413_/A2 _10137_/A _11788_/Q _06214_/C1 vssd1 vssd1 vccd1 vccd1
+ _06169_/X sky130_fd_sc_hd__o221a_1
XFILLER_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout720 _06459_/B1 vssd1 vssd1 vccd1 vccd1 _06630_/B1 sky130_fd_sc_hd__buf_4
Xfanout731 fanout738/X vssd1 vssd1 vccd1 vccd1 _06728_/B1 sky130_fd_sc_hd__buf_6
XFILLER_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout742 _06637_/A2 vssd1 vssd1 vccd1 vccd1 _06126_/B sky130_fd_sc_hd__buf_4
X_09928_ _11658_/Q _09770_/S _09890_/X _09927_/X vssd1 vssd1 vccd1 vccd1 _11658_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_104_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout753 _06214_/B1 vssd1 vssd1 vccd1 vccd1 _08994_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout764 _09132_/A vssd1 vssd1 vccd1 vccd1 _06739_/A2 sky130_fd_sc_hd__buf_4
Xfanout775 _09380_/A vssd1 vssd1 vccd1 vccd1 _06284_/B1 sky130_fd_sc_hd__buf_4
Xfanout786 _06806_/A2 vssd1 vssd1 vccd1 vccd1 _07540_/A sky130_fd_sc_hd__buf_6
X_09859_ _10713_/Q _09878_/A2 _09878_/B1 _10710_/Q vssd1 vssd1 vccd1 vccd1 _09859_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout797 _06641_/A2 vssd1 vssd1 vccd1 vccd1 _06152_/B sky130_fd_sc_hd__buf_6
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _09038_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_113 _09976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _08789_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _07010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_146 _05908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_157 _08840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11755_/CLK _11752_/D vssd1 vssd1 vccd1 vccd1 _11752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_168 input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_179 _10136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10773_/CLK _10703_/D vssd1 vssd1 vccd1 vccd1 _10703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11683_/CLK _11683_/D vssd1 vssd1 vccd1 vccd1 _11683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10634_ _11270_/CLK _10634_/D vssd1 vssd1 vccd1 vccd1 _10634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10565_ _11472_/CLK _10565_/D vssd1 vssd1 vccd1 vccd1 _10565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10496_ _11450_/CLK _10496_/D vssd1 vssd1 vccd1 vccd1 _10496_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_154_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ _11329_/CLK _11117_/D vssd1 vssd1 vccd1 vccd1 _11117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11048_ _11329_/CLK _11048_/D vssd1 vssd1 vccd1 vccd1 _11048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput8 ram_val_in[2] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_4
XFILLER_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05540_ _05630_/A2 _11352_/Q _11349_/Q _05079_/A _05538_/X vssd1 vssd1 vccd1 vccd1
+ _05543_/A sky130_fd_sc_hd__a221o_4
XFILLER_45_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05471_ _05471_/A _06942_/B _09679_/B vssd1 vssd1 vccd1 vccd1 _05472_/B sky130_fd_sc_hd__or3_1
XFILLER_75_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07210_ _10134_/A0 _07204_/B _07771_/B1 _10368_/Q vssd1 vssd1 vccd1 vccd1 _10368_/D
+ sky130_fd_sc_hd__a22o_1
X_08190_ _08193_/A _08190_/B vssd1 vssd1 vccd1 vccd1 _10929_/D sky130_fd_sc_hd__or2_1
XFILLER_20_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07141_ _07141_/A _07141_/B vssd1 vssd1 vccd1 vccd1 _07141_/X sky130_fd_sc_hd__and2_2
X_07072_ _10295_/Q _07078_/B vssd1 vssd1 vccd1 vccd1 _07072_/X sky130_fd_sc_hd__or2_1
XFILLER_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06023_ _11416_/Q _09132_/A vssd1 vssd1 vccd1 vccd1 _06023_/X sky130_fd_sc_hd__or2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07974_ _10810_/Q _07991_/S _07363_/S _07090_/A vssd1 vssd1 vccd1 vccd1 _10810_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09713_ _09713_/A _09713_/B _09713_/C _09713_/D vssd1 vssd1 vccd1 vccd1 _09721_/A
+ sky130_fd_sc_hd__or4_1
X_06925_ _10088_/A1 _10203_/Q _06934_/S vssd1 vssd1 vccd1 vccd1 _10203_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09644_ _10330_/Q _09573_/C _09570_/B _10326_/Q vssd1 vssd1 vccd1 vccd1 _09644_/X
+ sky130_fd_sc_hd__a22o_1
X_06856_ _10336_/Q _06856_/A2 _06710_/B _10803_/Q vssd1 vssd1 vccd1 vccd1 _06856_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05807_ _11061_/Q _06629_/A2 _06538_/B1 _10633_/Q _05806_/X vssd1 vssd1 vccd1 vccd1
+ _05807_/X sky130_fd_sc_hd__o221a_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09575_ _09576_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09908_/A sky130_fd_sc_hd__nor2_8
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06787_ _10529_/Q _06873_/A2 _06685_/B _11718_/Q _06786_/X vssd1 vssd1 vccd1 vccd1
+ _06787_/X sky130_fd_sc_hd__o221a_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08526_ _09101_/A1 _08529_/S _08525_/X _08947_/C1 vssd1 vssd1 vccd1 vccd1 _11112_/D
+ sky130_fd_sc_hd__o211a_1
X_05738_ _05749_/A _05751_/B _05745_/A vssd1 vssd1 vccd1 vccd1 _05738_/X sky130_fd_sc_hd__and3b_2
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08457_ _11078_/Q _07623_/X _07626_/S _07318_/B vssd1 vssd1 vccd1 vccd1 _11078_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05669_ _11204_/Q _05561_/Y _05585_/Y _11203_/Q vssd1 vssd1 vccd1 vccd1 _05669_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07408_ _10058_/A _07408_/B vssd1 vssd1 vccd1 vccd1 _10480_/D sky130_fd_sc_hd__or2_1
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08388_ _11035_/Q _08422_/B vssd1 vssd1 vccd1 vccd1 _08388_/X sky130_fd_sc_hd__or2_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07339_ _10435_/Q _07350_/S _07846_/S _07324_/B vssd1 vssd1 vccd1 vccd1 _10435_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_104_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10350_ _11457_/CLK _10350_/D vssd1 vssd1 vccd1 vccd1 _10350_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_136_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09009_ _11356_/Q _09013_/B vssd1 vssd1 vccd1 vccd1 _09009_/X sky130_fd_sc_hd__or2_1
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10281_ _10798_/CLK _10281_/D vssd1 vssd1 vccd1 vccd1 _10281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout550 _07790_/A vssd1 vssd1 vccd1 vccd1 _07926_/A sky130_fd_sc_hd__clkbuf_4
Xfanout561 fanout565/X vssd1 vssd1 vccd1 vccd1 _08771_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout572 _08670_/A vssd1 vssd1 vccd1 vccd1 _08781_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout583 _05818_/Y vssd1 vssd1 vccd1 vccd1 _06886_/A2 sky130_fd_sc_hd__buf_2
XFILLER_120_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout594 _07690_/Y vssd1 vssd1 vccd1 vccd1 _09038_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_101_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _11810_/CLK _11804_/D vssd1 vssd1 vccd1 vccd1 _11804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _11735_/CLK _11735_/D vssd1 vssd1 vccd1 vccd1 _11735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _11756_/CLK _11666_/D vssd1 vssd1 vccd1 vccd1 _11666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10617_ _11307_/CLK _10617_/D vssd1 vssd1 vccd1 vccd1 _10617_/Q sky130_fd_sc_hd__dfxtp_1
X_11597_ _11650_/CLK _11597_/D vssd1 vssd1 vccd1 vccd1 _11597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10548_ _10548_/CLK _10548_/D vssd1 vssd1 vccd1 vccd1 _10548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10479_ _11702_/CLK _10479_/D vssd1 vssd1 vccd1 vccd1 _10479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06710_ _10730_/Q _06710_/B vssd1 vssd1 vccd1 vccd1 _06710_/X sky130_fd_sc_hd__or2_1
XFILLER_77_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07690_ _07690_/A _07690_/B vssd1 vssd1 vccd1 vccd1 _07690_/Y sky130_fd_sc_hd__nand2_8
XFILLER_42_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06641_ _10934_/Q _06641_/A2 _08469_/B _11086_/Q _06640_/X vssd1 vssd1 vccd1 vccd1
+ _06641_/X sky130_fd_sc_hd__o221a_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _11538_/Q _09376_/B vssd1 vssd1 vccd1 vccd1 _09360_/X sky130_fd_sc_hd__or2_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06572_ _11202_/Q _06645_/A2 _09109_/A _11252_/Q vssd1 vssd1 vccd1 vccd1 _06572_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08311_ _08311_/A _10108_/B _10119_/C vssd1 vssd1 vccd1 vccd1 _08321_/S sky130_fd_sc_hd__or3_4
X_05523_ _05076_/A _11408_/Q _11403_/Q _05620_/B2 _05522_/X vssd1 vssd1 vccd1 vccd1
+ _05524_/B sky130_fd_sc_hd__a221o_4
X_09291_ _11497_/Q _09271_/X _09290_/X vssd1 vssd1 vccd1 vccd1 _11497_/D sky130_fd_sc_hd__a21o_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_13 _05968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05454_ _10767_/Q _09871_/A2 _09947_/B1 _10761_/Q vssd1 vssd1 vccd1 vccd1 _05454_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08242_ _08469_/A _08325_/B _08241_/Y _09267_/C1 vssd1 vssd1 vccd1 vccd1 _10954_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_24 _06883_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 _08683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_wb_clk_i clkbuf_leaf_88_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11243_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08173_ _07015_/A _10915_/Q _08181_/S vssd1 vssd1 vccd1 vccd1 _10915_/D sky130_fd_sc_hd__mux2_1
X_05385_ _10619_/Q _10618_/Q _05385_/S vssd1 vssd1 vccd1 vccd1 _05389_/A sky130_fd_sc_hd__mux2_1
XANTENNA_68 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 _11620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07124_ _10321_/Q _07126_/B _07186_/S _07333_/B vssd1 vssd1 vccd1 vccd1 _10321_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_107_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07055_ _10285_/Q _07047_/B _07490_/S _08811_/B2 vssd1 vssd1 vccd1 vccd1 _10285_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput120 _05644_/X vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_4
Xoutput131 _11611_/Q vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_4
Xoutput142 _11622_/Q vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__buf_4
X_06006_ _10584_/Q _06454_/A2 _06455_/B1 _10902_/Q vssd1 vssd1 vccd1 vccd1 _06006_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_115_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput153 _10218_/Q vssd1 vssd1 vccd1 vccd1 ram_val_out[0] sky130_fd_sc_hd__buf_4
XFILLER_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput164 _11584_/Q vssd1 vssd1 vccd1 vccd1 rom_addr[6] sky130_fd_sc_hd__buf_4
XFILLER_99_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput175 _11873_/X vssd1 vssd1 vccd1 vccd1 wb_rom_adrb[7] sky130_fd_sc_hd__buf_4
XFILLER_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput186 _05492_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_4
Xoutput197 _05502_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_4
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07957_ _07029_/X _10799_/Q _07961_/S vssd1 vssd1 vccd1 vccd1 _10799_/D sky130_fd_sc_hd__mux2_1
X_06908_ _10195_/Q _06922_/B vssd1 vssd1 vccd1 vccd1 _06908_/X sky130_fd_sc_hd__or2_1
X_07888_ _07932_/A1 _07890_/A2 _07887_/X _07932_/C1 vssd1 vssd1 vccd1 vccd1 _10762_/D
+ sky130_fd_sc_hd__o211a_1
X_09627_ _10802_/Q _09567_/A _09570_/A _10731_/Q vssd1 vssd1 vccd1 vccd1 _09627_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06839_ _06853_/A1 _10248_/Q _06853_/A3 _06838_/X _05819_/B vssd1 vssd1 vccd1 vccd1
+ _06839_/X sky130_fd_sc_hd__a32o_1
XFILLER_43_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09558_ _09558_/A _09600_/A vssd1 vssd1 vccd1 vccd1 _09827_/A sky130_fd_sc_hd__nand2_2
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08509_ _11104_/Q _08545_/B vssd1 vssd1 vccd1 vccd1 _08509_/X sky130_fd_sc_hd__or2_1
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09489_ _09525_/A _09489_/B _09489_/C vssd1 vssd1 vccd1 vccd1 _09490_/A sky130_fd_sc_hd__nand3_1
XFILLER_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11520_ _11527_/CLK _11520_/D vssd1 vssd1 vccd1 vccd1 _11520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ _11644_/CLK _11451_/D vssd1 vssd1 vccd1 vccd1 _11451_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10402_ _10808_/CLK _10402_/D vssd1 vssd1 vccd1 vccd1 _10402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11382_ _11428_/CLK _11382_/D vssd1 vssd1 vccd1 vccd1 _11382_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_152_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10333_ _10735_/CLK _10333_/D vssd1 vssd1 vccd1 vccd1 _10333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10264_ _11808_/CLK _10264_/D vssd1 vssd1 vccd1 vccd1 _10264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10195_ _11810_/CLK _10195_/D vssd1 vssd1 vccd1 vccd1 _10195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout380 _09214_/B vssd1 vssd1 vccd1 vccd1 _09226_/A sky130_fd_sc_hd__buf_6
Xfanout391 _08438_/A vssd1 vssd1 vccd1 vccd1 _08303_/A sky130_fd_sc_hd__buf_6
XFILLER_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11718_ _11719_/CLK _11718_/D vssd1 vssd1 vccd1 vccd1 _11718_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11649_ _11652_/CLK _11649_/D vssd1 vssd1 vccd1 vccd1 _11649_/Q sky130_fd_sc_hd__dfxtp_2
Xinput11 rom_value[10] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_2
Xinput22 rom_value[20] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput33 rom_value[30] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput44 wb_rom_val[11] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_2
X_05170_ _11184_/Q _11183_/Q _05326_/S vssd1 vssd1 vccd1 vccd1 _05176_/B sky130_fd_sc_hd__mux2_1
Xinput55 wb_rom_val[21] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput66 wb_rom_val[31] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_4
Xinput77 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__buf_6
Xinput88 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput99 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__buf_4
XFILLER_115_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08860_ _09276_/A1 _11287_/Q _08890_/S vssd1 vssd1 vccd1 vccd1 _08861_/B sky130_fd_sc_hd__mux2_1
XFILLER_112_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07811_ input101/X _10713_/Q _09200_/S vssd1 vssd1 vccd1 vccd1 _07812_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_106_wb_clk_i clkbuf_4_10__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11457_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08791_ _08933_/A1 _08792_/S _08790_/X _08791_/C1 vssd1 vssd1 vccd1 vccd1 _11251_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07742_ _10672_/Q _07760_/B vssd1 vssd1 vccd1 vccd1 _07742_/X sky130_fd_sc_hd__or2_1
XFILLER_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07673_ _08655_/B _08663_/S vssd1 vssd1 vccd1 vccd1 _07673_/Y sky130_fd_sc_hd__nor2_4
XFILLER_53_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09412_ _11333_/Q _11573_/Q _09414_/S vssd1 vssd1 vccd1 vccd1 _11573_/D sky130_fd_sc_hd__mux2_1
X_06624_ _11284_/Q _09359_/A _09977_/A _10843_/Q _06624_/C1 vssd1 vssd1 vccd1 vccd1
+ _06624_/X sky130_fd_sc_hd__o221a_1
XFILLER_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09343_ _11526_/Q _09343_/B vssd1 vssd1 vccd1 vccd1 _09343_/X sky130_fd_sc_hd__or2_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06555_ _11230_/Q _08650_/A _06640_/B1 _11142_/Q vssd1 vssd1 vccd1 vccd1 _06555_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05506_ _10251_/Q input63/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05506_/X sky130_fd_sc_hd__mux2_2
X_09274_ _11489_/Q _09288_/B vssd1 vssd1 vccd1 vccd1 _09274_/X sky130_fd_sc_hd__or2_1
X_06486_ _11044_/Q _09059_/A _08971_/A _10966_/Q vssd1 vssd1 vccd1 vccd1 _06486_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08225_ _08838_/A0 _10947_/Q _08225_/S vssd1 vssd1 vccd1 vccd1 _08226_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05437_ _10671_/Q _09883_/B1 _09950_/B1 _10662_/Q vssd1 vssd1 vccd1 vccd1 _05437_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05368_ _05368_/A _05368_/B vssd1 vssd1 vccd1 vccd1 _05368_/Y sky130_fd_sc_hd__nor2_8
X_08156_ _10904_/Q _08164_/B vssd1 vssd1 vccd1 vccd1 _08156_/X sky130_fd_sc_hd__or2_1
XFILLER_140_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07107_ _07107_/A _07107_/B vssd1 vssd1 vccd1 vccd1 _07335_/B sky130_fd_sc_hd__and2_4
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05299_ _11134_/Q _10450_/Q _06942_/A vssd1 vssd1 vccd1 vccd1 _05301_/C sky130_fd_sc_hd__mux2_1
X_08087_ _10869_/Q _08655_/B _08091_/C vssd1 vssd1 vccd1 vccd1 _08087_/X sky130_fd_sc_hd__or3_1
X_07038_ _10277_/Q _07037_/X _07038_/S vssd1 vssd1 vccd1 vccd1 _10277_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08989_ _11347_/Q _08989_/B vssd1 vssd1 vccd1 vccd1 _08989_/X sky130_fd_sc_hd__or2_1
XFILLER_29_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10951_ _11005_/CLK _10951_/D vssd1 vssd1 vccd1 vccd1 _10951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10882_ _10929_/CLK _10882_/D vssd1 vssd1 vccd1 vccd1 _10882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11503_ _11800_/CLK _11503_/D vssd1 vssd1 vccd1 vccd1 _11503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11434_ _11442_/CLK _11434_/D vssd1 vssd1 vccd1 vccd1 _11434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11365_ _11808_/CLK _11365_/D vssd1 vssd1 vccd1 vccd1 _11365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _10932_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10316_ _10735_/CLK _10316_/D vssd1 vssd1 vccd1 vccd1 _10316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11296_ _11325_/CLK _11296_/D vssd1 vssd1 vccd1 vccd1 _11296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10247_ _11474_/CLK _10247_/D vssd1 vssd1 vccd1 vccd1 _10247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10178_ _10178_/A1 _10176_/B _10178_/B1 vssd1 vssd1 vccd1 vccd1 _10178_/X sky130_fd_sc_hd__a21o_1
XFILLER_113_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06340_ _06663_/A _10230_/Q _06576_/A _06622_/A2 vssd1 vssd1 vccd1 vccd1 _06340_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06271_ _10649_/Q _06629_/A2 _06267_/X _06270_/X vssd1 vssd1 vccd1 vccd1 _06271_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08010_ _08833_/A _08010_/B vssd1 vssd1 vccd1 vccd1 _10829_/D sky130_fd_sc_hd__or2_1
X_05222_ _11054_/Q _11053_/Q _05427_/S vssd1 vssd1 vccd1 vccd1 _05223_/D sky130_fd_sc_hd__mux2_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05153_ _10946_/Q _10945_/Q _09680_/C vssd1 vssd1 vccd1 vccd1 _05156_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09961_ _11663_/Q _09820_/X _09963_/B vssd1 vssd1 vccd1 vccd1 _11663_/D sky130_fd_sc_hd__mux2_1
X_05084_ _05377_/S vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__clkinv_4
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08912_ _11315_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08912_/X sky130_fd_sc_hd__or2_1
XFILLER_48_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09892_ _11721_/Q _09567_/A _09948_/B1 _11709_/Q _09891_/X vssd1 vssd1 vccd1 vccd1
+ _09899_/A sky130_fd_sc_hd__a221o_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _09141_/A1 _08850_/S _08842_/X _08843_/C1 vssd1 vssd1 vccd1 vccd1 _11279_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08774_ _09141_/A1 _11243_/Q _08792_/S vssd1 vssd1 vccd1 vccd1 _08775_/B sky130_fd_sc_hd__mux2_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05986_ _11036_/Q _06696_/A2 _08245_/A _10958_/Q vssd1 vssd1 vccd1 vccd1 _05988_/B
+ sky130_fd_sc_hd__o22a_1
X_07725_ _08929_/A1 _07751_/A2 _07724_/X _09201_/A1 vssd1 vssd1 vccd1 vccd1 _10663_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07656_ _10620_/Q _07663_/S _07246_/S _07090_/A vssd1 vssd1 vccd1 vccd1 _10620_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11411_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06607_ _10290_/Q _09325_/A _09248_/A _10323_/Q vssd1 vssd1 vccd1 vccd1 _06607_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07587_ _07141_/A _10577_/Q _07589_/S vssd1 vssd1 vccd1 vccd1 _07588_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09326_ _09326_/A _10137_/B _10087_/C vssd1 vssd1 vccd1 vccd1 _09326_/X sky130_fd_sc_hd__or3_4
XFILLER_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06538_ _11068_/Q _06538_/A2 _06538_/B1 _11186_/Q vssd1 vssd1 vccd1 vccd1 _06538_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09257_ _11481_/Q _09249_/X _09256_/X vssd1 vssd1 vccd1 vccd1 _11481_/D sky130_fd_sc_hd__a21o_1
X_06469_ _10615_/Q _06641_/A2 _06639_/B1 _10454_/Q _06468_/X vssd1 vssd1 vccd1 vccd1
+ _06469_/X sky130_fd_sc_hd__o221a_1
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08208_ _08492_/A _08208_/B vssd1 vssd1 vccd1 vccd1 _10938_/D sky130_fd_sc_hd__or2_1
X_09188_ _07441_/A _09187_/X _09193_/A vssd1 vssd1 vccd1 vccd1 _11439_/D sky130_fd_sc_hd__o21a_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08139_ _08969_/A1 _08140_/S _08138_/X _08841_/C1 vssd1 vssd1 vccd1 vccd1 _10895_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11150_ _11151_/CLK _11150_/D vssd1 vssd1 vccd1 vccd1 _11150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10101_ _11752_/Q _10087_/X _10100_/X vssd1 vssd1 vccd1 vccd1 _11752_/D sky130_fd_sc_hd__a21o_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11081_ _11140_/CLK _11081_/D vssd1 vssd1 vccd1 vccd1 _11081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10032_ _11706_/Q _07061_/A _10051_/S vssd1 vssd1 vccd1 vccd1 _10033_/B sky130_fd_sc_hd__mux2_1
XFILLER_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10934_ _11584_/CLK _10934_/D vssd1 vssd1 vccd1 vccd1 _10934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10865_ _11485_/CLK _10865_/D vssd1 vssd1 vccd1 vccd1 _10865_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _11744_/CLK _10796_/D vssd1 vssd1 vccd1 vccd1 _10796_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11417_ _11792_/CLK _11417_/D vssd1 vssd1 vccd1 vccd1 _11417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11348_ _11497_/CLK _11348_/D vssd1 vssd1 vccd1 vccd1 _11348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11279_ _11280_/CLK _11279_/D vssd1 vssd1 vccd1 vccd1 _11279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05840_ _11803_/Q _10180_/A _05838_/X _05839_/X vssd1 vssd1 vccd1 vccd1 _05840_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05771_ _11802_/Q _10180_/A _05769_/X _05770_/X vssd1 vssd1 vccd1 vccd1 _05771_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07510_ _07916_/A _07510_/B vssd1 vssd1 vccd1 vccd1 _10539_/D sky130_fd_sc_hd__or2_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08490_ _09323_/A0 _08497_/S _08489_/X _09022_/C1 vssd1 vssd1 vccd1 vccd1 _11095_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07441_ _07441_/A _07537_/B vssd1 vssd1 vccd1 vccd1 _07441_/Y sky130_fd_sc_hd__nor2_4
XFILLER_22_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07372_ _10460_/Q _07309_/X _07373_/S vssd1 vssd1 vccd1 vccd1 _10460_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09111_ _09111_/A1 _09127_/B _08869_/A vssd1 vssd1 vccd1 vccd1 _09111_/X sky130_fd_sc_hd__a21o_1
X_06323_ _10941_/Q _06630_/A2 _06628_/B1 _11271_/Q vssd1 vssd1 vccd1 vccd1 _06323_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09042_ _09275_/A1 _09038_/X _09041_/X _09289_/C1 vssd1 vssd1 vccd1 vccd1 _11370_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06254_ _10845_/Q _06308_/A2 _10010_/A _11138_/Q _06253_/X vssd1 vssd1 vccd1 vccd1
+ _06255_/C sky130_fd_sc_hd__o221a_1
XFILLER_117_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05205_ _10902_/Q _10428_/Q _06939_/A vssd1 vssd1 vccd1 vccd1 _05205_/X sky130_fd_sc_hd__mux2_1
X_06185_ _11365_/Q _09016_/A _08994_/A _11355_/Q _06349_/C1 vssd1 vssd1 vccd1 vccd1
+ _06185_/X sky130_fd_sc_hd__o221a_1
XFILLER_132_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_121_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11477_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_05136_ _10644_/Q _10643_/Q _05413_/S vssd1 vssd1 vccd1 vccd1 _05140_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout902 _09081_/A vssd1 vssd1 vccd1 vccd1 _09358_/A sky130_fd_sc_hd__buf_12
X_09944_ _10371_/Q _09567_/B _09944_/B1 _10369_/Q _09941_/X vssd1 vssd1 vccd1 vccd1
+ _09957_/B sky130_fd_sc_hd__a221o_1
Xfanout913 _06297_/C1 vssd1 vssd1 vccd1 vccd1 _07151_/A sky130_fd_sc_hd__buf_6
Xfanout924 _06189_/A1 vssd1 vssd1 vccd1 vccd1 _06431_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout935 _07070_/A vssd1 vssd1 vccd1 vccd1 _08423_/A1 sky130_fd_sc_hd__buf_6
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout946 input94/X vssd1 vssd1 vccd1 vccd1 _08469_/A sky130_fd_sc_hd__buf_8
XFILLER_135_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout957 fanout958/X vssd1 vssd1 vccd1 vccd1 _09234_/A0 sky130_fd_sc_hd__buf_6
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09875_ _10556_/Q _09875_/A2 _09875_/B1 _10555_/Q _09874_/X vssd1 vssd1 vccd1 vccd1
+ _09880_/B sky130_fd_sc_hd__a221o_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout968 input90/X vssd1 vssd1 vccd1 vccd1 _07061_/A sky130_fd_sc_hd__buf_12
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout979 _08669_/A0 vssd1 vssd1 vccd1 vccd1 _07048_/A sky130_fd_sc_hd__buf_6
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08826_ _09323_/A0 _11271_/Q _08838_/S vssd1 vssd1 vccd1 vccd1 _08827_/B sky130_fd_sc_hd__mux2_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08757_ _08757_/A _08757_/B vssd1 vssd1 vccd1 vccd1 _11235_/D sky130_fd_sc_hd__or2_1
X_05969_ _11362_/Q _10087_/A _10137_/A _11352_/Q _06214_/C1 vssd1 vssd1 vccd1 vccd1
+ _05969_/X sky130_fd_sc_hd__o221a_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _10655_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07708_/X sky130_fd_sc_hd__or2_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08688_ _08875_/A _08688_/B vssd1 vssd1 vccd1 vccd1 _11198_/D sky130_fd_sc_hd__or2_1
XFILLER_57_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07639_ _08810_/A _08102_/S vssd1 vssd1 vccd1 vccd1 _07642_/S sky130_fd_sc_hd__nor2_8
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10650_ _11270_/CLK _10650_/D vssd1 vssd1 vccd1 vccd1 _10650_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09309_ _10175_/A1 _09293_/X _09308_/X _10175_/C1 vssd1 vssd1 vccd1 vccd1 _11505_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10581_ _11243_/CLK _10581_/D vssd1 vssd1 vccd1 vccd1 _10581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11202_ _11812_/CLK _11202_/D vssd1 vssd1 vccd1 vccd1 _11202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11133_ _11133_/CLK _11133_/D vssd1 vssd1 vccd1 vccd1 _11133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11064_ _11067_/CLK _11064_/D vssd1 vssd1 vccd1 vccd1 _11064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10015_ _10015_/A0 _11698_/Q _10028_/B vssd1 vssd1 vccd1 vccd1 _10016_/B sky130_fd_sc_hd__mux2_1
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10917_ _11779_/CLK _10917_/D vssd1 vssd1 vccd1 vccd1 _10917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10848_ _11308_/CLK _10848_/D vssd1 vssd1 vccd1 vccd1 _10848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10779_ _11457_/CLK _10779_/D vssd1 vssd1 vccd1 vccd1 _10779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07990_ _08193_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _10820_/D sky130_fd_sc_hd__or2_1
XFILLER_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06941_ _06941_/A _09431_/B _09679_/B _09681_/A vssd1 vssd1 vccd1 vccd1 _09538_/C
+ sky130_fd_sc_hd__and4_4
XFILLER_68_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09660_ _09650_/X _09659_/X _09959_/B vssd1 vssd1 vccd1 vccd1 _09660_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_95_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06872_ _10363_/Q _06872_/A2 _06685_/B _11745_/Q _06871_/X vssd1 vssd1 vccd1 vccd1
+ _06872_/X sky130_fd_sc_hd__o221a_1
XFILLER_68_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08611_ _09995_/A1 _11160_/Q _08621_/S vssd1 vssd1 vccd1 vccd1 _08612_/B sky130_fd_sc_hd__mux2_1
X_05823_ _11539_/Q _09359_/A _09293_/A _11499_/Q vssd1 vssd1 vccd1 vccd1 _05823_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09591_ _10510_/Q _09950_/B1 _09572_/D _10271_/Q vssd1 vssd1 vccd1 vccd1 _09593_/C
+ sky130_fd_sc_hd__a22o_1
X_08542_ _09237_/A0 _08537_/S _08541_/X _07003_/B vssd1 vssd1 vccd1 vccd1 _11120_/D
+ sky130_fd_sc_hd__o211a_1
X_05754_ _11792_/Q _10159_/A _06697_/B1 _11498_/Q vssd1 vssd1 vccd1 vccd1 _05754_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_70_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08473_ _11087_/Q _08503_/B vssd1 vssd1 vccd1 vccd1 _08473_/X sky130_fd_sc_hd__or2_1
X_05685_ _11158_/Q _05537_/Y _05633_/Y _11153_/Q vssd1 vssd1 vccd1 vccd1 _05685_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07424_ _10043_/A _07424_/B vssd1 vssd1 vccd1 vccd1 _10488_/D sky130_fd_sc_hd__or2_1
XFILLER_56_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07355_ _07102_/X _10448_/Q _07355_/S vssd1 vssd1 vccd1 vccd1 _10448_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06306_ _10622_/Q _06871_/A2 _06999_/A _10271_/Q vssd1 vssd1 vccd1 vccd1 _06309_/A
+ sky130_fd_sc_hd__o22a_1
X_07286_ _07930_/A _07286_/B vssd1 vssd1 vccd1 vccd1 _10411_/D sky130_fd_sc_hd__or2_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ _11363_/Q _09035_/B vssd1 vssd1 vccd1 vccd1 _09025_/X sky130_fd_sc_hd__or2_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06237_ _10354_/Q _06373_/B1 _07827_/A2 _10798_/Q _06236_/X vssd1 vssd1 vccd1 vccd1
+ _06237_/X sky130_fd_sc_hd__o221a_1
XFILLER_117_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06168_ _11524_/Q _09326_/A _06363_/A2 _11484_/Q vssd1 vssd1 vccd1 vccd1 _06168_/X
+ sky130_fd_sc_hd__o22a_1
X_05119_ _11175_/Q _10300_/Q _05380_/S vssd1 vssd1 vccd1 vccd1 _05123_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06099_ _11563_/Q _09391_/A _06284_/B1 _11553_/Q vssd1 vssd1 vccd1 vccd1 _06099_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout710 _10108_/C vssd1 vssd1 vccd1 vccd1 _10119_/C sky130_fd_sc_hd__buf_6
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout721 fanout726/X vssd1 vssd1 vccd1 vccd1 _06459_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_63_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout732 _06697_/B1 vssd1 vssd1 vccd1 vccd1 _06455_/B1 sky130_fd_sc_hd__buf_6
XFILLER_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09927_ _06948_/X _09908_/Y _09926_/Y vssd1 vssd1 vccd1 vccd1 _09927_/X sky130_fd_sc_hd__a21o_1
Xfanout743 _06640_/B1 vssd1 vssd1 vccd1 vccd1 _06637_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout754 fanout755/X vssd1 vssd1 vccd1 vccd1 _06214_/B1 sky130_fd_sc_hd__buf_4
Xfanout765 _05749_/X vssd1 vssd1 vccd1 vccd1 _09132_/A sky130_fd_sc_hd__buf_6
XFILLER_63_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout776 _08311_/A vssd1 vssd1 vccd1 vccd1 _09380_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout787 fanout793/X vssd1 vssd1 vccd1 vccd1 _06806_/A2 sky130_fd_sc_hd__buf_6
X_09858_ _11441_/Q _09877_/A2 _09877_/B1 _11442_/Q _09857_/X vssd1 vssd1 vccd1 vccd1
+ _09861_/C sky130_fd_sc_hd__a221o_1
XFILLER_111_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout798 _06998_/A vssd1 vssd1 vccd1 vccd1 _06731_/B1 sky130_fd_sc_hd__buf_6
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _11261_/Q _07015_/A _08820_/S vssd1 vssd1 vccd1 vccd1 _08810_/B sky130_fd_sc_hd__mux2_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09789_ _11649_/Q _09404_/Y _09788_/X _09681_/B vssd1 vssd1 vccd1 vccd1 _09789_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _09038_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 _06553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_125 _07059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_136 _07007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _05945_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11791_/CLK _11751_/D vssd1 vssd1 vccd1 vccd1 _11751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_158 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10702_ _10785_/CLK _10702_/D vssd1 vssd1 vccd1 vccd1 _10702_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11684_/CLK _11682_/D vssd1 vssd1 vccd1 vccd1 _11682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10633_ _10644_/CLK _10633_/D vssd1 vssd1 vccd1 vccd1 _10633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10564_ _11573_/CLK _10564_/D vssd1 vssd1 vccd1 vccd1 _10564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10495_ _11720_/CLK _10495_/D vssd1 vssd1 vccd1 vccd1 _10495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11116_ _11330_/CLK _11116_/D vssd1 vssd1 vccd1 vccd1 _11116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11047_ _11622_/CLK _11047_/D vssd1 vssd1 vccd1 vccd1 _11047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 ram_val_in[3] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_8
XFILLER_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05470_ _05470_/A _05470_/B vssd1 vssd1 vccd1 vccd1 _05474_/B sky130_fd_sc_hd__or2_4
XFILLER_33_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07140_ _10051_/A1 _07111_/X _07139_/X _07141_/B vssd1 vssd1 vccd1 vccd1 _10331_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07071_ _10294_/Q _07047_/B _07491_/S _07245_/B vssd1 vssd1 vccd1 vccd1 _10294_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_127_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06022_ _11680_/Q _08594_/A _06018_/X _06021_/X vssd1 vssd1 vccd1 vccd1 _06022_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07973_ _07143_/X _07901_/B _07972_/X vssd1 vssd1 vccd1 vccd1 _10809_/D sky130_fd_sc_hd__a21o_1
XFILLER_45_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ _10402_/Q _09567_/C _09872_/B1 _10399_/Q _09711_/X vssd1 vssd1 vccd1 vccd1
+ _09713_/D sky130_fd_sc_hd__a221o_1
X_06924_ _06924_/A _10108_/B _10180_/C vssd1 vssd1 vccd1 vccd1 _06934_/S sky130_fd_sc_hd__or3_4
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09643_ _10325_/Q _09565_/A _09571_/C _10331_/Q _09642_/X vssd1 vssd1 vccd1 vccd1
+ _09650_/A sky130_fd_sc_hd__a221o_2
XFILLER_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06855_ input74/X _06855_/B vssd1 vssd1 vccd1 vccd1 _06883_/C sky130_fd_sc_hd__nor2_8
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05806_ _10581_/Q _06454_/A2 _06539_/B1 _10591_/Q _06624_/C1 vssd1 vssd1 vccd1 vccd1
+ _05806_/X sky130_fd_sc_hd__o221a_2
X_09574_ _09574_/A _09574_/B _09574_/C _09574_/D vssd1 vssd1 vccd1 vccd1 _09576_/B
+ sky130_fd_sc_hd__or4_4
X_06786_ _10492_/Q _06872_/A2 _06856_/A2 _10332_/Q vssd1 vssd1 vccd1 vccd1 _06786_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08525_ _11112_/Q _08545_/B vssd1 vssd1 vccd1 vccd1 _08525_/X sky130_fd_sc_hd__or2_1
X_05737_ _05745_/A _05737_/B vssd1 vssd1 vccd1 vccd1 _05737_/X sky130_fd_sc_hd__or2_4
XFILLER_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08456_ _11077_/Q _08459_/S _07628_/S _07022_/B vssd1 vssd1 vccd1 vccd1 _11077_/D
+ sky130_fd_sc_hd__o22a_1
X_05668_ _05668_/A _05668_/B _05668_/C _05668_/D vssd1 vssd1 vccd1 vccd1 _05668_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07407_ _10021_/A0 _10480_/Q _07437_/S vssd1 vssd1 vccd1 vccd1 _07408_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08387_ _09114_/A1 _08404_/S _08386_/X _09092_/C1 vssd1 vssd1 vccd1 vccd1 _11034_/D
+ sky130_fd_sc_hd__o211a_1
X_05599_ _11684_/Q _05629_/A2 _05629_/B1 _11678_/Q vssd1 vssd1 vccd1 vccd1 _05599_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07338_ _08819_/A _07350_/S vssd1 vssd1 vccd1 vccd1 _07338_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07269_ _08929_/A1 _10403_/Q _07277_/S vssd1 vssd1 vccd1 vccd1 _07270_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09008_ _10150_/A1 _08994_/X _09007_/X _09032_/C1 vssd1 vssd1 vccd1 vccd1 _11355_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10280_ _11766_/CLK _10280_/D vssd1 vssd1 vccd1 vccd1 _10280_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout540 _10020_/A vssd1 vssd1 vccd1 vccd1 _10026_/A sky130_fd_sc_hd__buf_4
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout551 _07790_/A vssd1 vssd1 vccd1 vccd1 _07936_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout562 fanout565/X vssd1 vssd1 vccd1 vccd1 _08783_/A sky130_fd_sc_hd__buf_2
XFILLER_115_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout573 fanout578/X vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout584 _05818_/Y vssd1 vssd1 vccd1 vccd1 _06853_/A3 sky130_fd_sc_hd__buf_8
XFILLER_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout595 _07690_/Y vssd1 vssd1 vccd1 vccd1 _09271_/C sky130_fd_sc_hd__buf_4
XFILLER_58_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _11803_/CLK _11803_/D vssd1 vssd1 vccd1 vccd1 _11803_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11735_/CLK _11734_/D vssd1 vssd1 vccd1 vccd1 _11734_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _11665_/CLK _11665_/D vssd1 vssd1 vccd1 vccd1 _11665_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10616_ _11633_/CLK _10616_/D vssd1 vssd1 vccd1 vccd1 _10616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11596_ _11650_/CLK _11596_/D vssd1 vssd1 vccd1 vccd1 _11596_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10547_ _10782_/CLK _10547_/D vssd1 vssd1 vccd1 vccd1 _10547_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10478_ _11703_/CLK _10478_/D vssd1 vssd1 vccd1 vccd1 _10478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06640_ _11232_/Q _08650_/A _06640_/B1 _11144_/Q vssd1 vssd1 vccd1 vccd1 _06640_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06571_ _11326_/Q _06648_/A2 _10136_/A _11298_/Q _08243_/B vssd1 vssd1 vccd1 vccd1
+ _06571_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08310_ _10990_/Q _08301_/Y _08304_/Y _07019_/X vssd1 vssd1 vccd1 vccd1 _10990_/D
+ sky130_fd_sc_hd__a22o_1
X_05522_ _05619_/A1 _11411_/Q _11407_/Q _05619_/B2 _05520_/X vssd1 vssd1 vccd1 vccd1
+ _05522_/X sky130_fd_sc_hd__a221o_1
X_09290_ input117/X _09288_/B _09290_/B1 vssd1 vssd1 vccd1 vccd1 _09290_/X sky130_fd_sc_hd__a21o_1
XFILLER_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08241_ _08241_/A _08325_/B vssd1 vssd1 vccd1 vccd1 _08241_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_14 _06000_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05453_ _10809_/Q _09886_/B1 _09877_/B1 _10752_/Q vssd1 vssd1 vccd1 vccd1 _05453_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_25 _06883_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_36 _09692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_58 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ _07052_/A _10914_/Q _08182_/S vssd1 vssd1 vccd1 vccd1 _10914_/D sky130_fd_sc_hd__mux2_1
XANTENNA_69 _05644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05384_ _05384_/A _05384_/B _05384_/C _05384_/D vssd1 vssd1 vccd1 vccd1 _05390_/A
+ sky130_fd_sc_hd__or4_4
X_07123_ _10320_/Q _07135_/A2 _07123_/B1 _07318_/B vssd1 vssd1 vccd1 vccd1 _10320_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07054_ _10284_/Q _07078_/B _07496_/S _07095_/B vssd1 vssd1 vccd1 vccd1 _10284_/D
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_99_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _10765_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xoutput121 _05656_/X vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_4
XFILLER_115_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput132 _11612_/Q vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_4
X_06005_ _11090_/Q _06589_/A2 _06001_/X _06004_/X vssd1 vssd1 vccd1 vccd1 _06005_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput143 _11623_/Q vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_28_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11650_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xoutput154 _10219_/Q vssd1 vssd1 vccd1 vccd1 ram_val_out[1] sky130_fd_sc_hd__buf_4
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput165 _11585_/Q vssd1 vssd1 vccd1 vccd1 rom_addr[7] sky130_fd_sc_hd__buf_4
XFILLER_86_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput176 _11874_/X vssd1 vssd1 vccd1 vccd1 wb_rom_adrb[8] sky130_fd_sc_hd__buf_4
XFILLER_99_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput187 _05493_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_4
XFILLER_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput198 _05503_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_4
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07956_ _07019_/X _10798_/Q _07956_/S vssd1 vssd1 vccd1 vccd1 _10798_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06907_ _10182_/A0 _06903_/X _06906_/X _06990_/C1 vssd1 vssd1 vccd1 vccd1 _10194_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07887_ _10762_/Q _07901_/B vssd1 vssd1 vccd1 vccd1 _07887_/X sky130_fd_sc_hd__or2_1
XFILLER_56_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06838_ _06853_/A1 _10248_/Q _06852_/A3 _06743_/X _06837_/X vssd1 vssd1 vccd1 vccd1
+ _06838_/X sky130_fd_sc_hd__a32o_1
X_09626_ _09626_/A _09626_/B _09626_/C _09626_/D vssd1 vssd1 vccd1 vccd1 _09636_/A
+ sky130_fd_sc_hd__or4_1
X_09557_ _11646_/Q _11661_/Q vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__or2_1
X_06769_ _06853_/A1 _10243_/Q _06853_/A3 _06768_/X _05819_/B vssd1 vssd1 vccd1 vccd1
+ _06769_/X sky130_fd_sc_hd__a32o_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08508_ _08869_/A _08508_/B vssd1 vssd1 vccd1 vccd1 _11103_/D sky130_fd_sc_hd__or2_1
XFILLER_19_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09488_ _09553_/A _09668_/B _09488_/C _09959_/B vssd1 vssd1 vccd1 vccd1 _09488_/Y
+ sky130_fd_sc_hd__nor4_4
XFILLER_51_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08439_ _08439_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08439_/Y sky130_fd_sc_hd__nand2_2
XFILLER_12_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11450_ _11450_/CLK _11450_/D vssd1 vssd1 vccd1 vccd1 _11450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10401_ _11644_/CLK _10401_/D vssd1 vssd1 vccd1 vccd1 _10401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11381_ _11385_/CLK _11381_/D vssd1 vssd1 vccd1 vccd1 _11381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10332_ _11744_/CLK _10332_/D vssd1 vssd1 vccd1 vccd1 _10332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10263_ _11803_/CLK _10263_/D vssd1 vssd1 vccd1 vccd1 _10263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10194_ _11803_/CLK _10194_/D vssd1 vssd1 vccd1 vccd1 _10194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout370 _07012_/Y vssd1 vssd1 vccd1 vccd1 _08323_/A sky130_fd_sc_hd__buf_6
Xfanout381 _07613_/A vssd1 vssd1 vccd1 vccd1 _09214_/B sky130_fd_sc_hd__buf_8
Xfanout392 _07599_/A vssd1 vssd1 vccd1 vccd1 _08438_/A sky130_fd_sc_hd__buf_8
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11717_ _11720_/CLK _11717_/D vssd1 vssd1 vccd1 vccd1 _11717_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11648_ _11650_/CLK _11648_/D vssd1 vssd1 vccd1 vccd1 _11648_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput12 rom_value[11] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput23 rom_value[21] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
Xinput34 rom_value[31] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_2
Xinput45 wb_rom_val[12] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_2
X_11579_ _11652_/CLK _11579_/D vssd1 vssd1 vccd1 vccd1 _11579_/Q sky130_fd_sc_hd__dfxtp_2
Xinput56 wb_rom_val[22] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_4
Xinput67 wb_rom_val[3] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_2
XFILLER_155_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput78 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__buf_8
Xinput89 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_16
XFILLER_115_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07810_ _07930_/A _07810_/B vssd1 vssd1 vccd1 vccd1 _10712_/D sky130_fd_sc_hd__or2_1
X_08790_ _11251_/Q _08804_/B vssd1 vssd1 vccd1 vccd1 _08790_/X sky130_fd_sc_hd__or2_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07741_ _08893_/A1 _07751_/A2 _07740_/X _07884_/C1 vssd1 vssd1 vccd1 vccd1 _10671_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07672_ _09248_/A _08649_/C _10136_/C vssd1 vssd1 vccd1 vccd1 _08663_/S sky130_fd_sc_hd__and3_4
X_09411_ _09502_/A _11572_/Q _09414_/S vssd1 vssd1 vccd1 vccd1 _11572_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06623_ _11238_/Q _07300_/A _09249_/A _11188_/Q vssd1 vssd1 vccd1 vccd1 _06623_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09342_ _10175_/A1 _09326_/X _09341_/X _09993_/C1 vssd1 vssd1 vccd1 vccd1 _11525_/D
+ sky130_fd_sc_hd__o211a_1
X_06554_ _10932_/Q _06152_/B _06639_/B1 _10819_/Q _06553_/X vssd1 vssd1 vccd1 vccd1
+ _06554_/X sky130_fd_sc_hd__o221a_1
XFILLER_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05505_ _10250_/Q input62/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05505_/X sky130_fd_sc_hd__mux2_2
X_09273_ _11488_/Q _09271_/X _09272_/X vssd1 vssd1 vccd1 vccd1 _11488_/D sky130_fd_sc_hd__a21o_1
XFILLER_90_1349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06485_ _06479_/X _06484_/X input85/X vssd1 vssd1 vccd1 vccd1 _06485_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ _07107_/A _08225_/S _08223_/X _08351_/C1 vssd1 vssd1 vccd1 vccd1 _10946_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05436_ _10668_/Q _09944_/B1 _09872_/B1 _10658_/Q vssd1 vssd1 vccd1 vccd1 _05451_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08155_ _10171_/A1 _08162_/S _08154_/X _08843_/C1 vssd1 vssd1 vccd1 vccd1 _10903_/D
+ sky130_fd_sc_hd__o211a_1
X_05367_ _05367_/A _05367_/B _05367_/C _05367_/D vssd1 vssd1 vccd1 vccd1 _05368_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_140_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07106_ _10308_/Q _07105_/X _07109_/S vssd1 vssd1 vccd1 vccd1 _10308_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08086_ _08853_/A1 _08083_/S _08085_/X _09267_/C1 vssd1 vssd1 vccd1 vccd1 _10868_/D
+ sky130_fd_sc_hd__o211a_1
X_05298_ _10449_/Q _11133_/Q _06942_/B vssd1 vssd1 vccd1 vccd1 _05301_/B sky130_fd_sc_hd__mux2_1
XFILLER_134_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07037_ _09229_/A _07037_/B vssd1 vssd1 vccd1 vccd1 _07037_/X sky130_fd_sc_hd__and2_1
XFILLER_0_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08988_ _11346_/Q _08972_/X _08987_/X vssd1 vssd1 vccd1 vccd1 _11346_/D sky130_fd_sc_hd__a21o_1
XFILLER_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07939_ _07939_/A _08471_/B _10136_/C vssd1 vssd1 vccd1 vccd1 _08085_/B sky130_fd_sc_hd__and3_4
XFILLER_151_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10950_ _11234_/CLK _10950_/D vssd1 vssd1 vccd1 vccd1 _10950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ _10384_/Q _09571_/B _09572_/D _10622_/Q _09608_/X vssd1 vssd1 vccd1 vccd1
+ _09617_/C sky130_fd_sc_hd__a221o_1
X_10881_ _10929_/CLK _10881_/D vssd1 vssd1 vccd1 vccd1 _10881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11502_ _11801_/CLK _11502_/D vssd1 vssd1 vccd1 vccd1 _11502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11433_ _11473_/CLK _11433_/D vssd1 vssd1 vccd1 vccd1 _11433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11364_ _11808_/CLK _11364_/D vssd1 vssd1 vccd1 vccd1 _11364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10315_ _11703_/CLK _10315_/D vssd1 vssd1 vccd1 vccd1 _10315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11295_ _11325_/CLK _11295_/D vssd1 vssd1 vccd1 vccd1 _11295_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10246_ _11471_/CLK _10246_/D vssd1 vssd1 vccd1 vccd1 _10246_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10177_ _10177_/A1 _10159_/X _10176_/X _10177_/C1 vssd1 vssd1 vccd1 vccd1 _11800_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06270_ _11094_/Q _06629_/B1 _06268_/X _06269_/X vssd1 vssd1 vccd1 vccd1 _06270_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05221_ _11058_/Q _11057_/Q _11596_/Q vssd1 vssd1 vccd1 vccd1 _05223_/C sky130_fd_sc_hd__mux2_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05152_ _10936_/Q _10935_/Q _05427_/S vssd1 vssd1 vccd1 vccd1 _05156_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09960_ _11662_/Q _09817_/Y _09963_/B vssd1 vssd1 vccd1 vccd1 _11662_/D sky130_fd_sc_hd__mux2_1
X_05083_ _05430_/S vssd1 vssd1 vccd1 vccd1 _09679_/B sky130_fd_sc_hd__inv_6
X_08911_ _09275_/A1 _08945_/A2 _08910_/X _09092_/C1 vssd1 vssd1 vccd1 vccd1 _11314_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09891_ _11743_/Q _09566_/C _09573_/C _11716_/Q vssd1 vssd1 vccd1 vccd1 _09891_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _11279_/Q _08852_/B vssd1 vssd1 vccd1 vccd1 _08842_/X sky130_fd_sc_hd__or2_1
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08773_/A _08773_/B vssd1 vssd1 vccd1 vccd1 _11242_/D sky130_fd_sc_hd__or2_1
X_05985_ _11316_/Q _08907_/A _08855_/A _11288_/Q _06718_/C1 vssd1 vssd1 vccd1 vccd1
+ _05988_/A sky130_fd_sc_hd__o221a_1
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07724_ _10663_/Q _07760_/B vssd1 vssd1 vccd1 vccd1 _07724_/X sky130_fd_sc_hd__or2_1
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ _08901_/A1 _10619_/Q _07655_/S vssd1 vssd1 vccd1 vccd1 _10619_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06606_ _11468_/Q _06649_/A2 _06602_/X _06605_/X vssd1 vssd1 vccd1 vccd1 _06606_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07586_ _07934_/A _07586_/B vssd1 vssd1 vccd1 vccd1 _10576_/D sky130_fd_sc_hd__or2_1
XFILLER_0_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09325_ _09325_/A _10136_/B _10158_/C vssd1 vssd1 vccd1 vccd1 _09343_/B sky130_fd_sc_hd__and3_4
XFILLER_94_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06537_ _11612_/Q _06622_/A2 _06535_/B _06622_/B2 _06536_/X vssd1 vssd1 vccd1 vccd1
+ _10234_/D sky130_fd_sc_hd__a221o_1
XFILLER_142_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09256_ _09256_/A1 _09266_/B _10150_/B1 vssd1 vssd1 vccd1 vccd1 _09256_/X sky130_fd_sc_hd__a21o_1
X_06468_ _10609_/Q _06468_/B vssd1 vssd1 vccd1 vccd1 _06468_/X sky130_fd_sc_hd__or2_1
XFILLER_103_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08207_ _10112_/A0 _10938_/Q _08225_/S vssd1 vssd1 vccd1 vccd1 _08208_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11810_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_05419_ _11236_/Q _11235_/Q _05419_/S vssd1 vssd1 vccd1 vccd1 _05422_/B sky130_fd_sc_hd__mux2_1
X_09187_ _07143_/A _11439_/Q _09187_/S vssd1 vssd1 vccd1 vccd1 _09187_/X sky130_fd_sc_hd__mux2_1
X_06399_ _10443_/Q _06634_/B1 _06731_/B1 _10597_/Q _06550_/C1 vssd1 vssd1 vccd1 vccd1
+ _06399_/X sky130_fd_sc_hd__o221a_1
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08138_ _10895_/Q _08637_/C vssd1 vssd1 vccd1 vccd1 _08138_/X sky130_fd_sc_hd__or2_1
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08069_ _10860_/Q _08426_/B vssd1 vssd1 vccd1 vccd1 _08069_/X sky130_fd_sc_hd__or2_1
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10100_ _10150_/A1 _10104_/B _10156_/B1 vssd1 vssd1 vccd1 vccd1 _10100_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11080_ _11781_/CLK _11080_/D vssd1 vssd1 vccd1 vccd1 _11080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10031_ _10039_/A _10031_/B vssd1 vssd1 vccd1 vccd1 _11705_/D sky130_fd_sc_hd__or2_1
XFILLER_114_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10933_ _11584_/CLK _10933_/D vssd1 vssd1 vccd1 vccd1 _10933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10864_ _11234_/CLK _10864_/D vssd1 vssd1 vccd1 vccd1 _10864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10795_ _10798_/CLK _10795_/D vssd1 vssd1 vccd1 vccd1 _10795_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11416_ _11792_/CLK _11416_/D vssd1 vssd1 vccd1 vccd1 _11416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11347_ _11497_/CLK _11347_/D vssd1 vssd1 vccd1 vccd1 _11347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11278_ _11601_/CLK _11278_/D vssd1 vssd1 vccd1 vccd1 _11278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10229_ _10981_/CLK _10229_/D vssd1 vssd1 vccd1 vccd1 _10229_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__buf_2
XFILLER_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05770_ _10256_/Q _06230_/A2 _06903_/A _10193_/Q vssd1 vssd1 vccd1 vccd1 _05770_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07440_ _07440_/A _07854_/B vssd1 vssd1 vccd1 vccd1 _07440_/X sky130_fd_sc_hd__or2_1
XFILLER_62_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07371_ _10459_/Q _07229_/X _07373_/S vssd1 vssd1 vccd1 vccd1 _10459_/D sky130_fd_sc_hd__mux2_1
X_09110_ _09110_/A _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09110_/X sky130_fd_sc_hd__or3_4
XFILLER_148_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06322_ _11063_/Q _06538_/A2 _06318_/X _06321_/X vssd1 vssd1 vccd1 vccd1 _06322_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09041_ _11370_/Q _09055_/B vssd1 vssd1 vccd1 vccd1 _09041_/X sky130_fd_sc_hd__or2_1
X_06253_ _10467_/Q _06371_/A2 _07827_/A2 _10982_/Q vssd1 vssd1 vccd1 vccd1 _06253_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05204_ _05199_/X _05204_/B _05204_/C _05204_/D vssd1 vssd1 vccd1 vccd1 _05204_/X
+ sky130_fd_sc_hd__and4b_4
X_06184_ _11564_/Q _09391_/A _06284_/B1 _11554_/Q vssd1 vssd1 vccd1 vccd1 _06184_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05135_ _05135_/A _05135_/B vssd1 vssd1 vccd1 vccd1 _05135_/Y sky130_fd_sc_hd__nor2_8
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09943_ _10695_/Q _09572_/B _09566_/D _10376_/Q _09942_/X vssd1 vssd1 vccd1 vccd1
+ _09957_/A sky130_fd_sc_hd__a221o_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout903 _09081_/A vssd1 vssd1 vccd1 vccd1 _06646_/A2 sky130_fd_sc_hd__clkbuf_16
Xfanout914 _06265_/C1 vssd1 vssd1 vccd1 vccd1 _06349_/C1 sky130_fd_sc_hd__buf_4
XFILLER_98_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout925 _06189_/A1 vssd1 vssd1 vccd1 vccd1 _07690_/A sky130_fd_sc_hd__buf_12
Xfanout936 _07070_/A vssd1 vssd1 vccd1 vccd1 _08947_/A1 sky130_fd_sc_hd__buf_2
XFILLER_86_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _10554_/Q _09874_/A2 _09567_/C _10563_/Q vssd1 vssd1 vccd1 vccd1 _09874_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout947 input94/X vssd1 vssd1 vccd1 vccd1 _08665_/A sky130_fd_sc_hd__buf_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout958 input93/X vssd1 vssd1 vccd1 vccd1 fanout958/X sky130_fd_sc_hd__buf_12
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout969 input90/X vssd1 vssd1 vccd1 vccd1 _08970_/A1 sky130_fd_sc_hd__buf_4
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08825_ _09971_/A0 _08838_/S _08824_/X _08831_/C1 vssd1 vssd1 vccd1 vccd1 _11270_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05968_ _11561_/Q _09391_/A _06284_/B1 _11551_/Q vssd1 vssd1 vccd1 vccd1 _05968_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_45_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08756_ _07104_/A _11235_/Q _08760_/S vssd1 vssd1 vccd1 vccd1 _08757_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07707_ _07303_/A _07751_/A2 _07706_/X _07894_/C1 vssd1 vssd1 vccd1 vccd1 _10654_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05899_ _11688_/Q _09998_/A _06924_/A _11735_/Q _06344_/C1 vssd1 vssd1 vccd1 vccd1
+ _05899_/X sky130_fd_sc_hd__o221a_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _09101_/A1 _11198_/Q _08707_/S vssd1 vssd1 vccd1 vccd1 _08688_/B sky130_fd_sc_hd__mux2_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07638_ _09358_/A _08649_/B _08560_/C vssd1 vssd1 vccd1 vccd1 _07638_/X sky130_fd_sc_hd__and3_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07569_ _09182_/A0 _10568_/Q _07591_/S vssd1 vssd1 vccd1 vccd1 _07570_/B sky130_fd_sc_hd__mux2_1
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09308_ _11505_/Q _09310_/B vssd1 vssd1 vccd1 vccd1 _09308_/X sky130_fd_sc_hd__or2_1
X_10580_ _11458_/CLK _10580_/D vssd1 vssd1 vccd1 vccd1 _10580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09239_ _07243_/B _07172_/S _09227_/Y _11471_/Q _09229_/A vssd1 vssd1 vccd1 vccd1
+ _11471_/D sky130_fd_sc_hd__o221a_1
XFILLER_103_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11201_ _11251_/CLK _11201_/D vssd1 vssd1 vccd1 vccd1 _11201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11132_ _11177_/CLK _11132_/D vssd1 vssd1 vccd1 vccd1 _11132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11063_ _11067_/CLK _11063_/D vssd1 vssd1 vccd1 vccd1 _11063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10014_ _10026_/A _10014_/B vssd1 vssd1 vccd1 vccd1 _11697_/D sky130_fd_sc_hd__or2_1
XFILLER_77_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10916_ _11781_/CLK _10916_/D vssd1 vssd1 vccd1 vccd1 _10916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10847_ _11140_/CLK _10847_/D vssd1 vssd1 vccd1 vccd1 _10847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10778_ _10782_/CLK _10778_/D vssd1 vssd1 vccd1 vccd1 _10778_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_73_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06940_ _09538_/A _08956_/B vssd1 vssd1 vccd1 vccd1 _09553_/A sky130_fd_sc_hd__nand2_4
XFILLER_140_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06871_ _10632_/Q _06871_/A2 _06871_/B1 _10737_/Q vssd1 vssd1 vccd1 vccd1 _06871_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_95_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05822_ _06450_/A _10223_/Q vssd1 vssd1 vccd1 vccd1 _05822_/X sky130_fd_sc_hd__and2_1
X_08610_ _08987_/A1 _08623_/S _08609_/X _08937_/C1 vssd1 vssd1 vccd1 vccd1 _11159_/D
+ sky130_fd_sc_hd__o211a_1
X_09590_ _10514_/Q _09568_/C _09565_/B _10513_/Q _09589_/X vssd1 vssd1 vccd1 vccd1
+ _09593_/B sky130_fd_sc_hd__a221o_1
XFILLER_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05753_ _11746_/Q _10087_/A _06214_/B1 _11782_/Q _06214_/C1 vssd1 vssd1 vccd1 vccd1
+ _05753_/X sky130_fd_sc_hd__o221a_1
X_08541_ _11120_/Q _08545_/B vssd1 vssd1 vccd1 vccd1 _08541_/X sky130_fd_sc_hd__or2_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08472_ _08472_/A _08665_/C _09038_/C vssd1 vssd1 vccd1 vccd1 _08472_/X sky130_fd_sc_hd__or3_2
XFILLER_63_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05684_ _11160_/Q _05549_/Y _05603_/Y _11156_/Q _05683_/X vssd1 vssd1 vccd1 vccd1
+ _05692_/B sky130_fd_sc_hd__a221o_1
XFILLER_1_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07423_ _07028_/A _10488_/Q _07437_/S vssd1 vssd1 vccd1 vccd1 _07424_/B sky130_fd_sc_hd__mux2_1
XFILLER_17_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07354_ _09232_/B2 _10447_/Q _07355_/S vssd1 vssd1 vccd1 vccd1 _10447_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06305_ _10365_/Q _06370_/A2 _07827_/A2 _10721_/Q vssd1 vssd1 vccd1 vccd1 _06305_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07285_ _10047_/A1 _10411_/Q _09184_/S vssd1 vssd1 vccd1 vccd1 _07286_/B sky130_fd_sc_hd__mux2_1
XFILLER_104_1348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09024_ _09256_/A1 _09016_/X _09023_/X _09267_/C1 vssd1 vssd1 vccd1 vccd1 _11362_/D
+ sky130_fd_sc_hd__o211a_1
X_06236_ _10270_/Q _06999_/A _06857_/B1 _11702_/Q vssd1 vssd1 vccd1 vccd1 _06236_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06167_ _11029_/Q _06538_/A2 _06163_/X _06166_/X vssd1 vssd1 vccd1 vccd1 _06167_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05118_ _05118_/A _05118_/B _05118_/C _05118_/D vssd1 vssd1 vccd1 vccd1 _05124_/A
+ sky130_fd_sc_hd__or4_4
X_06098_ _11513_/Q _09314_/A _06094_/X _06097_/X vssd1 vssd1 vccd1 vccd1 _06098_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_137_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout700 _05427_/S vssd1 vssd1 vccd1 vccd1 _05391_/S sky130_fd_sc_hd__clkbuf_16
Xfanout711 _05787_/X vssd1 vssd1 vccd1 vccd1 _07082_/A sky130_fd_sc_hd__buf_8
Xfanout722 _08097_/A vssd1 vssd1 vccd1 vccd1 _09347_/A sky130_fd_sc_hd__clkbuf_8
X_09926_ _09908_/A _09925_/X _09770_/S vssd1 vssd1 vccd1 vccd1 _09926_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout733 _06697_/B1 vssd1 vssd1 vccd1 vccd1 _09293_/A sky130_fd_sc_hd__buf_6
Xfanout744 fanout755/X vssd1 vssd1 vccd1 vccd1 _06640_/B1 sky130_fd_sc_hd__buf_6
Xfanout755 _05749_/X vssd1 vssd1 vccd1 vccd1 fanout755/X sky130_fd_sc_hd__buf_8
XFILLER_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout766 _10136_/A vssd1 vssd1 vccd1 vccd1 _08560_/A sky130_fd_sc_hd__buf_12
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout777 _08300_/A vssd1 vssd1 vccd1 vccd1 _08311_/A sky130_fd_sc_hd__buf_4
XFILLER_24_1338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _10716_/Q _09876_/A2 _09876_/B1 _10705_/Q vssd1 vssd1 vccd1 vccd1 _09857_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout788 _08245_/A vssd1 vssd1 vccd1 vccd1 _06363_/A2 sky130_fd_sc_hd__buf_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout799 _06641_/A2 vssd1 vssd1 vccd1 vccd1 _06998_/A sky130_fd_sc_hd__buf_6
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _11260_/Q _08820_/S _07630_/Y _07617_/B vssd1 vssd1 vccd1 vccd1 _11260_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09788_ _11650_/Q _09771_/Y _09787_/X _09554_/B _09406_/B vssd1 vssd1 vccd1 vccd1
+ _09788_/X sky130_fd_sc_hd__o221a_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _07057_/A _08748_/S _08738_/X _08578_/A vssd1 vssd1 vccd1 vccd1 _11226_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _05413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_115 _06553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _07298_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_137 _10142_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _05962_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11791_/CLK _11750_/D vssd1 vssd1 vccd1 vccd1 _11750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_159 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _11575_/CLK _10701_/D vssd1 vssd1 vccd1 vccd1 _10701_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11681_ _11684_/CLK _11681_/D vssd1 vssd1 vccd1 vccd1 _11681_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10632_ _11711_/CLK _10632_/D vssd1 vssd1 vccd1 vccd1 _10632_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10563_ _11573_/CLK _10563_/D vssd1 vssd1 vccd1 vccd1 _10563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _11720_/CLK _10494_/D vssd1 vssd1 vccd1 vccd1 _10494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11115_ _11330_/CLK _11115_/D vssd1 vssd1 vccd1 vccd1 _11115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11046_ _11812_/CLK _11046_/D vssd1 vssd1 vccd1 vccd1 _11046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ _07070_/A _07107_/B vssd1 vssd1 vccd1 vccd1 _07245_/B sky130_fd_sc_hd__and2_1
XFILLER_69_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06021_ _11542_/Q _06219_/A2 _06019_/X _06020_/X vssd1 vssd1 vccd1 vccd1 _06021_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07972_ _10809_/Q _09227_/A _07966_/S _09228_/A vssd1 vssd1 vccd1 vccd1 _07972_/X
+ sky130_fd_sc_hd__a31o_1
X_09711_ _10414_/Q _09879_/A2 _09878_/A2 _11437_/Q vssd1 vssd1 vccd1 vccd1 _09711_/X
+ sky130_fd_sc_hd__a22o_1
X_06923_ _10106_/A1 _06903_/X _06922_/X _06996_/C1 vssd1 vssd1 vccd1 vccd1 _10202_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09642_ _10336_/Q _09909_/A2 _09572_/B _10332_/Q vssd1 vssd1 vccd1 vccd1 _09642_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06854_ _11657_/Q _06704_/B _06853_/X vssd1 vssd1 vccd1 vccd1 _10249_/D sky130_fd_sc_hd__a21o_1
XFILLER_82_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05805_ _10417_/Q _06541_/A2 _06589_/A2 _10949_/Q _05804_/X vssd1 vssd1 vccd1 vccd1
+ _05805_/X sky130_fd_sc_hd__o221a_1
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06785_ _10695_/Q _07203_/A _06858_/B1 _10519_/Q vssd1 vssd1 vccd1 vccd1 _06785_/X
+ sky130_fd_sc_hd__o22a_1
X_09573_ _09573_/A _09573_/B _09573_/C _09573_/D vssd1 vssd1 vccd1 vccd1 _09574_/D
+ sky130_fd_sc_hd__or4_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08524_ _08783_/A _08524_/B vssd1 vssd1 vccd1 vccd1 _11111_/D sky130_fd_sc_hd__or2_1
X_05736_ _05745_/A _05737_/B vssd1 vssd1 vccd1 vccd1 _05736_/Y sky130_fd_sc_hd__nor2_8
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08455_ _11076_/Q _08459_/S _07628_/S _08811_/B2 vssd1 vssd1 vccd1 vccd1 _11076_/D
+ sky130_fd_sc_hd__o22a_1
X_05667_ _11245_/Q _05537_/Y _05573_/Y _11248_/Q _05666_/X vssd1 vssd1 vccd1 vccd1
+ _05668_/D sky130_fd_sc_hd__a221o_2
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07406_ _07476_/A _07406_/B vssd1 vssd1 vccd1 vccd1 _10479_/D sky130_fd_sc_hd__or2_1
X_08386_ _11034_/Q _08422_/B vssd1 vssd1 vccd1 vccd1 _08386_/X sky130_fd_sc_hd__or2_1
XFILLER_149_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05598_ _11683_/Q _05628_/A2 _05628_/B1 _11680_/Q vssd1 vssd1 vccd1 vccd1 _05598_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07337_ _09358_/A _08560_/C _07847_/C vssd1 vssd1 vccd1 vccd1 _07337_/X sky130_fd_sc_hd__and3_4
XFILLER_13_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07268_ _07796_/A _07268_/B vssd1 vssd1 vccd1 vccd1 _10402_/D sky130_fd_sc_hd__or2_1
XFILLER_87_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06219_ _11396_/Q _06219_/A2 _09132_/A _11419_/Q vssd1 vssd1 vccd1 vccd1 _06219_/X
+ sky130_fd_sc_hd__o22a_1
X_09007_ _11355_/Q _09013_/B vssd1 vssd1 vccd1 vccd1 _09007_/X sky130_fd_sc_hd__or2_1
XFILLER_151_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07199_ _07147_/A _07191_/B _07192_/A _10361_/Q _07451_/A vssd1 vssd1 vccd1 vccd1
+ _10361_/D sky130_fd_sc_hd__a221o_1
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout530 fanout536/X vssd1 vssd1 vccd1 vccd1 _08492_/A sky130_fd_sc_hd__buf_4
XFILLER_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout541 _10020_/A vssd1 vssd1 vccd1 vccd1 _07928_/A sky130_fd_sc_hd__buf_4
XFILLER_115_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09909_ _10362_/Q _09909_/A2 _09944_/B1 _10358_/Q vssd1 vssd1 vccd1 vccd1 _09909_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout552 _07818_/A vssd1 vssd1 vccd1 vccd1 _07796_/A sky130_fd_sc_hd__clkbuf_4
Xfanout563 fanout565/X vssd1 vssd1 vccd1 vccd1 _10166_/B1 sky130_fd_sc_hd__buf_4
XFILLER_28_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout574 fanout578/X vssd1 vssd1 vccd1 vccd1 _08873_/A sky130_fd_sc_hd__buf_4
XFILLER_24_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout585 _05818_/Y vssd1 vssd1 vccd1 vccd1 _06622_/B2 sky130_fd_sc_hd__buf_4
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout596 _07689_/Y vssd1 vssd1 vccd1 vccd1 _09037_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_24_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_9__f_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_9__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _11809_/CLK _11802_/D vssd1 vssd1 vccd1 vccd1 _11802_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _11733_/CLK _11733_/D vssd1 vssd1 vccd1 vccd1 _11733_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11664_ _11665_/CLK _11664_/D vssd1 vssd1 vccd1 vccd1 _11664_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10615_ _10932_/CLK _10615_/D vssd1 vssd1 vccd1 vccd1 _10615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11595_ _11601_/CLK _11595_/D vssd1 vssd1 vccd1 vccd1 _11595_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10546_ _11457_/CLK _10546_/D vssd1 vssd1 vccd1 vccd1 _10546_/Q sky130_fd_sc_hd__dfxtp_1
X_10477_ _11706_/CLK _10477_/D vssd1 vssd1 vccd1 vccd1 _10477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11029_ _11067_/CLK _11029_/D vssd1 vssd1 vccd1 vccd1 _11029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06570_ _11046_/Q _05736_/Y _05746_/X _10968_/Q vssd1 vssd1 vccd1 vccd1 _06570_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05521_ _05618_/A1 _11405_/Q _11402_/Q _05606_/B2 _05519_/X vssd1 vssd1 vccd1 vccd1
+ _05524_/A sky130_fd_sc_hd__a221o_4
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08240_ _08761_/A _08240_/B vssd1 vssd1 vccd1 vccd1 _10953_/D sky130_fd_sc_hd__or2_1
X_05452_ _05452_/A _05452_/B vssd1 vssd1 vccd1 vccd1 _05474_/A sky130_fd_sc_hd__or2_4
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_15 _06151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _10159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_37 _09811_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ _07092_/A _10913_/Q _08181_/S vssd1 vssd1 vccd1 vccd1 _10913_/D sky130_fd_sc_hd__mux2_1
XANTENNA_48 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05383_ _10469_/Q _10468_/Q _05432_/S vssd1 vssd1 vccd1 vccd1 _05384_/D sky130_fd_sc_hd__mux2_2
XANTENNA_59 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07122_ _10319_/Q _07126_/B _07186_/S _07316_/B vssd1 vssd1 vccd1 vccd1 _10319_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07053_ _10283_/Q _07078_/B _07496_/S _07617_/B vssd1 vssd1 vccd1 vccd1 _10283_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput122 _05668_/X vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_4
X_06004_ _11146_/Q _07692_/A _06002_/X _06003_/X vssd1 vssd1 vccd1 vccd1 _06004_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput133 _11613_/Q vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_4
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput144 _11587_/Q vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__buf_4
XFILLER_138_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput155 _10220_/Q vssd1 vssd1 vccd1 vccd1 ram_val_out[2] sky130_fd_sc_hd__buf_4
XFILLER_99_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput166 _11586_/Q vssd1 vssd1 vccd1 vccd1 rom_addr[8] sky130_fd_sc_hd__buf_4
Xoutput177 _06890_/Y vssd1 vssd1 vccd1 vccd1 wb_rom_csb sky130_fd_sc_hd__buf_4
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput188 _05494_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_4
XFILLER_138_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput199 _05504_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_4
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_68_wb_clk_i clkbuf_leaf_69_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11431_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07955_ _07309_/X _10797_/Q _07956_/S vssd1 vssd1 vccd1 vccd1 _10797_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06906_ _10194_/Q _06922_/B vssd1 vssd1 vccd1 vccd1 _06906_/X sky130_fd_sc_hd__or2_1
XFILLER_96_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07886_ _08423_/A1 _07966_/S _07885_/X _07932_/C1 vssd1 vssd1 vccd1 vccd1 _10761_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09625_ _10798_/Q _09571_/B _09572_/D _10721_/Q vssd1 vssd1 vccd1 vccd1 _09626_/D
+ sky130_fd_sc_hd__a22o_1
X_06837_ _06832_/X _06833_/X _06836_/X _06831_/X vssd1 vssd1 vccd1 vccd1 _06837_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09556_ _11646_/Q _11661_/Q vssd1 vssd1 vccd1 vccd1 _09558_/A sky130_fd_sc_hd__nand2_1
X_06768_ _06853_/A1 _10243_/Q _06852_/A3 _06743_/X _06767_/X vssd1 vssd1 vccd1 vccd1
+ _06768_/X sky130_fd_sc_hd__a32o_1
XFILLER_145_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08507_ _09111_/A1 _11103_/Q _08529_/S vssd1 vssd1 vccd1 vccd1 _08508_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05719_ _10971_/Q _05579_/Y _05597_/Y _10962_/Q vssd1 vssd1 vccd1 vccd1 _05719_/X
+ sky130_fd_sc_hd__a22o_1
X_09487_ _09522_/B _09522_/C vssd1 vssd1 vccd1 vccd1 _09489_/B sky130_fd_sc_hd__nor2_1
X_06699_ _11206_/Q _06736_/A2 _06735_/B1 _11169_/Q _06698_/X vssd1 vssd1 vccd1 vccd1
+ _06699_/X sky130_fd_sc_hd__o221a_1
XFILLER_145_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08438_ _08438_/A _08438_/B vssd1 vssd1 vccd1 vccd1 _08438_/Y sky130_fd_sc_hd__nor2_2
XFILLER_145_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08369_ _08757_/A _08369_/B vssd1 vssd1 vccd1 vccd1 _11026_/D sky130_fd_sc_hd__or2_1
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ _10773_/CLK _10400_/D vssd1 vssd1 vccd1 vccd1 _10400_/Q sky130_fd_sc_hd__dfxtp_2
X_11380_ _11385_/CLK _11380_/D vssd1 vssd1 vccd1 vccd1 _11380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10331_ _11719_/CLK _10331_/D vssd1 vssd1 vccd1 vccd1 _10331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ _11803_/CLK _10262_/D vssd1 vssd1 vccd1 vccd1 _10262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10193_ _11755_/CLK _10193_/D vssd1 vssd1 vccd1 vccd1 _10193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout360 _09270_/B vssd1 vssd1 vccd1 vccd1 _10136_/B sky130_fd_sc_hd__buf_8
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout371 _09227_/A vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__buf_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout382 _07011_/Y vssd1 vssd1 vccd1 vccd1 _07613_/A sky130_fd_sc_hd__buf_6
Xfanout393 _09228_/A vssd1 vssd1 vccd1 vccd1 _07451_/A sky130_fd_sc_hd__buf_6
XFILLER_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11716_/CLK _11716_/D vssd1 vssd1 vccd1 vccd1 _11716_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11647_ _11650_/CLK _11647_/D vssd1 vssd1 vccd1 vccd1 _11647_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_11_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput13 rom_value[12] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput24 rom_value[22] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput35 rom_value[3] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput46 wb_rom_val[13] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_4
X_11578_ _11652_/CLK _11578_/D vssd1 vssd1 vccd1 vccd1 _11578_/Q sky130_fd_sc_hd__dfxtp_2
Xinput57 wb_rom_val[23] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput68 wb_rom_val[4] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_2
XFILLER_156_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10529_ _11722_/CLK _10529_/D vssd1 vssd1 vccd1 vccd1 _10529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput79 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__buf_2
XFILLER_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07740_ _10671_/Q _07750_/B vssd1 vssd1 vccd1 vccd1 _07740_/X sky130_fd_sc_hd__or2_1
XFILLER_42_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07671_ _10632_/Q _07665_/S _07249_/S _07043_/B vssd1 vssd1 vccd1 vccd1 _10632_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09410_ _09511_/C _11571_/Q _09414_/S vssd1 vssd1 vccd1 vccd1 _11571_/D sky130_fd_sc_hd__mux2_1
XFILLER_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06622_ _11614_/Q _06622_/A2 _06620_/X _06622_/B2 _06621_/X vssd1 vssd1 vccd1 vccd1
+ _10236_/D sky130_fd_sc_hd__a221o_1
XFILLER_20_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09341_ _11525_/Q _09343_/B vssd1 vssd1 vccd1 vccd1 _09341_/X sky130_fd_sc_hd__or2_1
X_06553_ _10885_/Q _06553_/B vssd1 vssd1 vccd1 vccd1 _06553_/X sky130_fd_sc_hd__or2_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05504_ _10249_/Q input61/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05504_/X sky130_fd_sc_hd__mux2_2
XFILLER_139_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09272_ _10161_/A1 _09288_/B _09290_/B1 vssd1 vssd1 vccd1 vccd1 _09272_/X sky130_fd_sc_hd__a21o_1
X_06484_ _11706_/Q _08560_/A _06480_/X _06483_/X vssd1 vssd1 vccd1 vccd1 _06484_/X
+ sky130_fd_sc_hd__a211o_2
Xclkbuf_leaf_115_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11719_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05435_ _10663_/Q _09573_/B _09571_/C _10675_/Q vssd1 vssd1 vccd1 vccd1 _05435_/X
+ sky130_fd_sc_hd__a22o_1
X_08223_ _10946_/Q _08902_/C vssd1 vssd1 vccd1 vccd1 _08223_/X sky130_fd_sc_hd__or2_1
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05366_ _11272_/Q _11271_/Q _05432_/S vssd1 vssd1 vccd1 vccd1 _05367_/D sky130_fd_sc_hd__mux2_1
X_08154_ _10903_/Q _08164_/B vssd1 vssd1 vccd1 vccd1 _08154_/X sky130_fd_sc_hd__or2_1
XFILLER_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07105_ _07318_/A _07333_/B vssd1 vssd1 vccd1 vccd1 _07105_/X sky130_fd_sc_hd__or2_4
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08085_ _10868_/Q _08085_/B vssd1 vssd1 vccd1 vccd1 _08085_/X sky130_fd_sc_hd__or2_1
XFILLER_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05297_ _11124_/Q _11123_/Q _05380_/S vssd1 vssd1 vccd1 vccd1 _05301_/A sky130_fd_sc_hd__mux2_1
X_07036_ _07036_/A _10056_/A vssd1 vssd1 vccd1 vccd1 _07037_/B sky130_fd_sc_hd__or2_4
XFILLER_134_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08987_ _08987_/A1 _08989_/B _09129_/B1 vssd1 vssd1 vccd1 vccd1 _08987_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07938_ _10056_/A _07938_/B vssd1 vssd1 vccd1 vccd1 _10786_/D sky130_fd_sc_hd__or2_1
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07869_ _10753_/Q _07883_/B vssd1 vssd1 vccd1 vccd1 _07869_/X sky130_fd_sc_hd__or2_1
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09608_ _10629_/Q _09571_/A _09950_/B1 _10623_/Q vssd1 vssd1 vccd1 vccd1 _09608_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10880_ _10932_/CLK _10880_/D vssd1 vssd1 vccd1 vccd1 _10880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09539_ _09539_/A _09539_/B _09668_/B _09668_/D vssd1 vssd1 vccd1 vccd1 _09539_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_52_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ _11801_/CLK _11501_/D vssd1 vssd1 vccd1 vccd1 _11501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11432_ _11473_/CLK _11432_/D vssd1 vssd1 vccd1 vccd1 _11432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11363_ _11366_/CLK _11363_/D vssd1 vssd1 vccd1 vccd1 _11363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10314_ _10812_/CLK _10314_/D vssd1 vssd1 vccd1 vccd1 _10314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11294_ _11319_/CLK _11294_/D vssd1 vssd1 vccd1 vccd1 _11294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10245_ _11474_/CLK _10245_/D vssd1 vssd1 vccd1 vccd1 _10245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10176_ _11800_/Q _10176_/B vssd1 vssd1 vccd1 vccd1 _10176_/X sky130_fd_sc_hd__or2_1
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05220_ _05085_/Y _11060_/Q _10859_/Q _09430_/B vssd1 vssd1 vccd1 vccd1 _05224_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05151_ _05151_/A _05151_/B _05151_/C _05151_/D vssd1 vssd1 vccd1 vccd1 _05157_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_155_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05082_ _09680_/C vssd1 vssd1 vccd1 vccd1 _09431_/B sky130_fd_sc_hd__clkinv_4
XFILLER_131_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08910_ _11314_/Q _08946_/B vssd1 vssd1 vccd1 vccd1 _08910_/X sky130_fd_sc_hd__or2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _11662_/Q _09851_/Y _09889_/Y input6/X _09870_/Y vssd1 vssd1 vccd1 vccd1
+ _09890_/X sky130_fd_sc_hd__a221o_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08469_/A _08838_/S _08840_/X _08841_/C1 vssd1 vssd1 vccd1 vccd1 _11278_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _09090_/A1 _11242_/Q _08792_/S vssd1 vssd1 vccd1 vccd1 _08773_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05984_ _05976_/X _05977_/X _05978_/X _05983_/X vssd1 vssd1 vccd1 vccd1 _05984_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07723_ _09129_/A1 _07751_/A2 _07722_/X _07884_/C1 vssd1 vssd1 vccd1 vccd1 _10662_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07654_ _07100_/X _10618_/Q _07655_/S vssd1 vssd1 vccd1 vccd1 _10618_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06605_ _10756_/Q _06648_/A2 _06604_/X _06873_/D1 vssd1 vssd1 vccd1 vccd1 _06605_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07585_ _07933_/A0 _10576_/Q _07591_/S vssd1 vssd1 vccd1 vccd1 _07586_/B sky130_fd_sc_hd__mux2_1
XFILLER_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09324_ _10118_/A0 _11517_/Q _09324_/S vssd1 vssd1 vccd1 vccd1 _11517_/D sky130_fd_sc_hd__mux2_1
X_06536_ _06576_/A _06533_/X _06535_/X _06664_/C1 vssd1 vssd1 vccd1 vccd1 _06536_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09255_ _09364_/A1 _09249_/X _09254_/X _10155_/C1 vssd1 vssd1 vccd1 vccd1 _11480_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06467_ _06467_/A _06467_/B _06467_/C vssd1 vssd1 vccd1 vccd1 _06467_/X sky130_fd_sc_hd__and3_1
XFILLER_142_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08206_ _08579_/A0 _08225_/S _08205_/X _09022_/C1 vssd1 vssd1 vccd1 vccd1 _10937_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05418_ _10418_/Q _10417_/Q _05418_/S vssd1 vssd1 vccd1 vccd1 _05422_/A sky130_fd_sc_hd__mux2_1
X_06398_ _10918_/Q _06591_/A2 _05865_/B _11775_/Q vssd1 vssd1 vccd1 vccd1 _06398_/X
+ sky130_fd_sc_hd__o22a_1
X_09186_ _07187_/B _09175_/B _09175_/Y _11438_/Q _09228_/A vssd1 vssd1 vccd1 vccd1
+ _11438_/D sky130_fd_sc_hd__a221o_1
XFILLER_105_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05349_ _11142_/Q _11141_/Q _05349_/S vssd1 vssd1 vccd1 vccd1 _05356_/A sky130_fd_sc_hd__mux2_1
X_08137_ _10190_/A0 _08140_/S _08136_/X _08841_/C1 vssd1 vssd1 vccd1 vccd1 _10894_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_wb_clk_i clkbuf_leaf_85_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11622_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08068_ _08833_/A _08068_/B vssd1 vssd1 vccd1 vccd1 _10859_/D sky130_fd_sc_hd__or2_1
XFILLER_134_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11136_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07019_ _08303_/A _07232_/B vssd1 vssd1 vccd1 vccd1 _07019_/X sky130_fd_sc_hd__or2_4
XFILLER_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10030_ _11705_/Q _07059_/A _10051_/S vssd1 vssd1 vccd1 vccd1 _10031_/B sky130_fd_sc_hd__mux2_1
XFILLER_66_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10932_ _10932_/CLK _10932_/D vssd1 vssd1 vccd1 vccd1 _10932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10863_ _11284_/CLK _10863_/D vssd1 vssd1 vccd1 vccd1 _10863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _11235_/CLK _10794_/D vssd1 vssd1 vccd1 vccd1 _10794_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11415_ _11792_/CLK _11415_/D vssd1 vssd1 vccd1 vccd1 _11415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11346_ _11495_/CLK _11346_/D vssd1 vssd1 vccd1 vccd1 _11346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11277_ _11601_/CLK _11277_/D vssd1 vssd1 vccd1 vccd1 _11277_/Q sky130_fd_sc_hd__dfxtp_1
X_10228_ _11233_/CLK _10228_/D vssd1 vssd1 vccd1 vccd1 _10228_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10159_ _10159_/A _10159_/B _10159_/C vssd1 vssd1 vccd1 vccd1 _10159_/X sky130_fd_sc_hd__or3_4
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07370_ _10458_/Q _07227_/X _07373_/S vssd1 vssd1 vccd1 vccd1 _10458_/D sky130_fd_sc_hd__mux2_1
X_06321_ _11005_/Q _06504_/B1 _06319_/X _06320_/X vssd1 vssd1 vccd1 vccd1 _06321_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09040_ _11369_/Q _09038_/X _09039_/X vssd1 vssd1 vccd1 vccd1 _11369_/D sky130_fd_sc_hd__a21o_1
X_06252_ _10880_/Q _06513_/A2 _06636_/A2 _10928_/Q _07083_/B vssd1 vssd1 vccd1 vccd1
+ _06255_/B sky130_fd_sc_hd__o221a_1
XFILLER_148_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05203_ _05203_/A _05203_/B vssd1 vssd1 vccd1 vccd1 _05204_/D sky130_fd_sc_hd__nor2_1
XFILLER_141_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06183_ _11514_/Q _08472_/A _06179_/X _06182_/X vssd1 vssd1 vccd1 vccd1 _06183_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_102_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05134_ _05134_/A _05134_/B _05134_/C _05134_/D vssd1 vssd1 vccd1 vccd1 _05135_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_89_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09942_ _10683_/Q _09566_/B _09571_/D _10686_/Q vssd1 vssd1 vccd1 vccd1 _09942_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout904 _05738_/X vssd1 vssd1 vccd1 vccd1 _09081_/A sky130_fd_sc_hd__buf_12
Xfanout915 _06265_/C1 vssd1 vssd1 vccd1 vccd1 _06214_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout926 _05091_/Y vssd1 vssd1 vccd1 vccd1 _06189_/A1 sky130_fd_sc_hd__buf_12
XFILLER_131_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout937 input98/X vssd1 vssd1 vccd1 vccd1 _07070_/A sky130_fd_sc_hd__buf_12
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09873_ _10558_/Q _09873_/A2 _09873_/B1 _10567_/Q _09872_/X vssd1 vssd1 vccd1 vccd1
+ _09880_/A sky130_fd_sc_hd__a221o_1
XFILLER_98_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout948 _08939_/A1 vssd1 vssd1 vccd1 vccd1 _07211_/A sky130_fd_sc_hd__buf_6
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout959 _08661_/A vssd1 vssd1 vccd1 vccd1 _07107_/A sky130_fd_sc_hd__buf_8
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _11270_/Q _08840_/B vssd1 vssd1 vccd1 vccd1 _08824_/X sky130_fd_sc_hd__or2_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08755_ _08757_/A _08755_/B vssd1 vssd1 vccd1 vccd1 _11234_/D sky130_fd_sc_hd__or2_1
XFILLER_85_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05967_ _11511_/Q _09314_/A _05963_/X _05966_/X vssd1 vssd1 vccd1 vccd1 _05967_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07706_ _10654_/Q _07750_/B vssd1 vssd1 vccd1 vccd1 _07706_/X sky130_fd_sc_hd__or2_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_130_wb_clk_i clkbuf_4_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11766_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08686_ _08771_/A _08686_/B vssd1 vssd1 vccd1 vccd1 _11197_/D sky130_fd_sc_hd__or2_1
X_05898_ _11725_/Q _08200_/A _09347_/A _11530_/Q vssd1 vssd1 vccd1 vccd1 _05898_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_57_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _10606_/Q _08901_/A1 _07637_/S vssd1 vssd1 vccd1 vccd1 _10606_/D sky130_fd_sc_hd__mux2_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07568_ _08536_/A _07568_/B vssd1 vssd1 vccd1 vccd1 _10567_/D sky130_fd_sc_hd__or2_1
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09307_ _11504_/Q _09293_/X _09306_/X vssd1 vssd1 vccd1 vccd1 _11504_/D sky130_fd_sc_hd__a21o_1
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06519_ _11443_/Q _09059_/A _09109_/A _10541_/Q _06518_/X vssd1 vssd1 vccd1 vccd1
+ _06519_/X sky130_fd_sc_hd__a221o_1
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07499_ _10534_/Q _07537_/B vssd1 vssd1 vccd1 vccd1 _07499_/X sky130_fd_sc_hd__or2_1
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09238_ _07441_/A _09237_/X _09241_/B1 vssd1 vssd1 vccd1 vccd1 _11470_/D sky130_fd_sc_hd__o21a_1
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ _10175_/A1 _09171_/B _10166_/B1 vssd1 vssd1 vccd1 vccd1 _09169_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11200_ _11683_/CLK _11200_/D vssd1 vssd1 vccd1 vccd1 _11200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11131_ _11780_/CLK _11131_/D vssd1 vssd1 vccd1 vccd1 _11131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11062_ _11067_/CLK _11062_/D vssd1 vssd1 vccd1 vccd1 _11062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10013_ _10013_/A0 _11697_/Q _10028_/B vssd1 vssd1 vccd1 vccd1 _10014_/B sky130_fd_sc_hd__mux2_1
XFILLER_95_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ _11770_/CLK _10915_/D vssd1 vssd1 vccd1 vccd1 _10915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10846_ _11310_/CLK _10846_/D vssd1 vssd1 vccd1 vccd1 _10846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ _11661_/CLK _10777_/D vssd1 vssd1 vccd1 vccd1 _10777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11329_ _11329_/CLK _11329_/D vssd1 vssd1 vccd1 vccd1 _11329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06870_ _10378_/Q _07904_/A _06870_/B1 _10279_/Q _06869_/X vssd1 vssd1 vccd1 vccd1
+ _06870_/X sky130_fd_sc_hd__o221a_1
XFILLER_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05821_ _05731_/X _06886_/A2 _06622_/A2 _05644_/X _05817_/X vssd1 vssd1 vccd1 vccd1
+ _10222_/D sky130_fd_sc_hd__a221o_1
XFILLER_83_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08540_ _09216_/A0 _08529_/S _08539_/X _08921_/C1 vssd1 vssd1 vccd1 vccd1 _11119_/D
+ sky130_fd_sc_hd__o211a_1
X_05752_ _11518_/Q _09326_/A _06363_/A2 _11478_/Q vssd1 vssd1 vccd1 vccd1 _05752_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08471_ _08560_/A _08471_/B _09037_/C vssd1 vssd1 vccd1 vccd1 _08503_/B sky130_fd_sc_hd__and3_4
X_05683_ _11167_/Q _05561_/Y _05567_/Y _11155_/Q vssd1 vssd1 vccd1 vccd1 _05683_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07422_ _10043_/A _07422_/B vssd1 vssd1 vccd1 vccd1 _10487_/D sky130_fd_sc_hd__or2_1
XFILLER_50_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07353_ _07664_/A _07353_/B vssd1 vssd1 vccd1 vccd1 _07353_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06304_ _11442_/Q _07778_/A _06303_/X _06808_/C1 vssd1 vssd1 vccd1 vccd1 _06304_/X
+ sky130_fd_sc_hd__o211a_1
X_07284_ _07926_/A _07284_/B vssd1 vssd1 vccd1 vccd1 _10410_/D sky130_fd_sc_hd__or2_1
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09023_ _11362_/Q _09035_/B vssd1 vssd1 vccd1 vccd1 _09023_/X sky130_fd_sc_hd__or2_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06235_ _10688_/Q _06370_/A2 _06371_/A2 _10384_/Q vssd1 vssd1 vccd1 vccd1 _06235_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06166_ _10594_/Q _06166_/A2 _06165_/X _06265_/C1 vssd1 vssd1 vccd1 vccd1 _06166_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05117_ _11177_/Q _10302_/Q _05393_/S vssd1 vssd1 vccd1 vccd1 _05118_/D sky130_fd_sc_hd__mux2_1
X_06097_ _11761_/Q _10108_/A _06095_/X _06096_/X vssd1 vssd1 vccd1 vccd1 _06097_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout701 _11594_/Q vssd1 vssd1 vccd1 vccd1 _05427_/S sky130_fd_sc_hd__buf_12
XFILLER_137_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09925_ _09925_/A _09925_/B _09925_/C _09925_/D vssd1 vssd1 vccd1 vccd1 _09925_/X
+ sky130_fd_sc_hd__or4_4
Xfanout712 _07081_/A vssd1 vssd1 vccd1 vccd1 _06619_/A1 sky130_fd_sc_hd__buf_4
XFILLER_131_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout723 fanout726/X vssd1 vssd1 vccd1 vccd1 _08097_/A sky130_fd_sc_hd__buf_4
XFILLER_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout734 fanout738/X vssd1 vssd1 vccd1 vccd1 _06697_/B1 sky130_fd_sc_hd__buf_6
Xfanout745 fanout755/X vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__buf_8
XFILLER_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout756 _06857_/B1 vssd1 vssd1 vccd1 vccd1 _06685_/B sky130_fd_sc_hd__buf_6
Xfanout767 _10136_/A vssd1 vssd1 vccd1 vccd1 _09131_/A sky130_fd_sc_hd__clkbuf_16
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _10699_/Q _09875_/A2 _09875_/B1 _10698_/Q _09855_/X vssd1 vssd1 vccd1 vccd1
+ _09861_/B sky130_fd_sc_hd__a221o_1
Xfanout778 fanout782/X vssd1 vssd1 vccd1 vccd1 _08300_/A sky130_fd_sc_hd__buf_4
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout789 fanout793/X vssd1 vssd1 vccd1 vccd1 _08245_/A sky130_fd_sc_hd__buf_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08807_ _08819_/A _08807_/B vssd1 vssd1 vccd1 vccd1 _11259_/D sky130_fd_sc_hd__or2_1
XFILLER_74_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8__f_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_8__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09787_ _05426_/S _09672_/B _09674_/A _11591_/Q vssd1 vssd1 vccd1 vccd1 _09787_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06999_ _06999_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _07483_/S sky130_fd_sc_hd__or2_4
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08738_ _11226_/Q _08750_/B vssd1 vssd1 vccd1 vccd1 _08738_/X sky130_fd_sc_hd__or2_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_105 _05413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_116 _06194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _09214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _05135_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _06075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ _08669_/A0 _11189_/Q _08707_/S vssd1 vssd1 vccd1 vccd1 _08670_/B sky130_fd_sc_hd__mux2_1
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _11471_/CLK _10700_/D vssd1 vssd1 vccd1 vccd1 _10700_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11683_/CLK _11680_/D vssd1 vssd1 vccd1 vccd1 _11680_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10631_ _11474_/CLK _10631_/D vssd1 vssd1 vccd1 vccd1 _10631_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10562_ _11622_/CLK _10562_/D vssd1 vssd1 vccd1 vccd1 _10562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10493_ _11719_/CLK _10493_/D vssd1 vssd1 vccd1 vccd1 _10493_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11114_ _11428_/CLK _11114_/D vssd1 vssd1 vccd1 vccd1 _11114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11045_ _11243_/CLK _11045_/D vssd1 vssd1 vccd1 vccd1 _11045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10829_ _11632_/CLK _10829_/D vssd1 vssd1 vccd1 vccd1 _10829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06020_ _11796_/Q _09154_/A _09293_/A _11502_/Q vssd1 vssd1 vccd1 vccd1 _06020_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_154_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07971_ _07441_/A _07970_/X _09241_/B1 vssd1 vssd1 vccd1 vccd1 _10808_/D sky130_fd_sc_hd__o21a_1
XFILLER_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09710_ _10411_/Q _09879_/B1 _09878_/B1 _10408_/Q _09709_/X vssd1 vssd1 vccd1 vccd1
+ _09713_/C sky130_fd_sc_hd__a221o_1
X_06922_ _10202_/Q _06922_/B vssd1 vssd1 vccd1 vccd1 _06922_/X sky130_fd_sc_hd__or2_1
XFILLER_68_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09641_ _09599_/X _09618_/X _09640_/X vssd1 vssd1 vccd1 vccd1 _09641_/Y sky130_fd_sc_hd__a21oi_2
X_06853_ _06853_/A1 _10249_/Q _06853_/A3 _06852_/X _05819_/B vssd1 vssd1 vccd1 vccd1
+ _06853_/X sky130_fd_sc_hd__a32o_1
XFILLER_28_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05804_ _10861_/Q _06540_/A2 _06540_/B1 _10427_/Q vssd1 vssd1 vccd1 vccd1 _05804_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_23_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09572_ _09572_/A _09572_/B _09572_/C _09572_/D vssd1 vssd1 vccd1 vccd1 _09574_/C
+ sky130_fd_sc_hd__or4_1
X_06784_ _11622_/Q _06704_/B _06783_/X vssd1 vssd1 vccd1 vccd1 _10244_/D sky130_fd_sc_hd__a21o_1
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08523_ _09172_/A1 _11111_/Q _08537_/S vssd1 vssd1 vccd1 vccd1 _08524_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05735_ _05749_/A _05751_/B vssd1 vssd1 vccd1 vccd1 _05737_/B sky130_fd_sc_hd__nand2_4
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08454_ _11075_/Q _08459_/S _07628_/S _07095_/B vssd1 vssd1 vccd1 vccd1 _11075_/D
+ sky130_fd_sc_hd__o22a_1
X_05666_ _11258_/Q _05518_/Y _05524_/Y _11249_/Q vssd1 vssd1 vccd1 vccd1 _05666_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07405_ _07052_/A _10479_/Q _07429_/S vssd1 vssd1 vccd1 vccd1 _07406_/B sky130_fd_sc_hd__mux2_1
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08385_ _08941_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _11033_/D sky130_fd_sc_hd__or2_1
X_05597_ _05597_/A _05597_/B vssd1 vssd1 vccd1 vccd1 _05597_/Y sky130_fd_sc_hd__nor2_8
XFILLER_52_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07336_ _10434_/Q _07323_/Y _07325_/Y _07335_/X vssd1 vssd1 vccd1 vccd1 _10434_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07267_ _09129_/A1 _10402_/Q _07277_/S vssd1 vssd1 vccd1 vccd1 _07268_/B sky130_fd_sc_hd__mux2_1
X_09006_ _10149_/A1 _08994_/X _09005_/X _09036_/C1 vssd1 vssd1 vccd1 vccd1 _11354_/D
+ sky130_fd_sc_hd__o211a_1
X_06218_ _11386_/Q _08383_/A vssd1 vssd1 vccd1 vccd1 _06218_/X sky130_fd_sc_hd__or2_1
X_07198_ _10051_/A1 _07191_/B _07192_/A _10360_/Q _07451_/A vssd1 vssd1 vccd1 vccd1
+ _10360_/D sky130_fd_sc_hd__a221o_1
XFILLER_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06149_ _10466_/Q _06371_/A2 _07827_/A2 _10981_/Q vssd1 vssd1 vccd1 vccd1 _06149_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout520 _07420_/A vssd1 vssd1 vccd1 vccd1 _10050_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout531 _10150_/B1 vssd1 vssd1 vccd1 vccd1 _08761_/A sky130_fd_sc_hd__buf_4
XFILLER_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout542 _10020_/A vssd1 vssd1 vccd1 vccd1 _07920_/A sky130_fd_sc_hd__clkbuf_2
X_09908_ _09908_/A _09908_/B vssd1 vssd1 vccd1 vccd1 _09908_/Y sky130_fd_sc_hd__nor2_2
Xfanout553 _07790_/A vssd1 vssd1 vccd1 vccd1 _07818_/A sky130_fd_sc_hd__buf_2
Xfanout564 fanout565/X vssd1 vssd1 vccd1 vccd1 _09173_/B1 sky130_fd_sc_hd__buf_2
XFILLER_24_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout575 fanout578/X vssd1 vssd1 vccd1 vccd1 _09290_/B1 sky130_fd_sc_hd__buf_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout586 _05734_/X vssd1 vssd1 vccd1 vccd1 _05816_/A sky130_fd_sc_hd__clkbuf_8
Xfanout597 _07689_/Y vssd1 vssd1 vccd1 vccd1 _09270_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_111_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09839_ _11461_/Q _09871_/A2 _09567_/C _10773_/Q _09838_/X vssd1 vssd1 vccd1 vccd1
+ _09842_/C sky130_fd_sc_hd__a221o_1
XFILLER_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _11801_/CLK _11801_/D vssd1 vssd1 vccd1 vccd1 _11801_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11733_/CLK _11732_/D vssd1 vssd1 vccd1 vccd1 _11732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11663_/CLK _11663_/D vssd1 vssd1 vccd1 vccd1 _11663_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10614_ _11310_/CLK _10614_/D vssd1 vssd1 vccd1 vccd1 _10614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11594_ _11650_/CLK _11594_/D vssd1 vssd1 vccd1 vccd1 _11594_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_70_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10545_ _10773_/CLK _10545_/D vssd1 vssd1 vccd1 vccd1 _10545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10476_ _11661_/CLK _10476_/D vssd1 vssd1 vccd1 vccd1 _10476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11028_ _11067_/CLK _11028_/D vssd1 vssd1 vccd1 vccd1 _11028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05520_ _09552_/A1 _11410_/Q _11404_/Q _05078_/A vssd1 vssd1 vccd1 vccd1 _05520_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05451_ _05451_/A _05451_/B _05451_/C _05451_/D vssd1 vssd1 vccd1 vccd1 _05452_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_75_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_16 _06200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_27 _07008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ _07010_/A _10912_/Q _08181_/S vssd1 vssd1 vccd1 vccd1 _10912_/D sky130_fd_sc_hd__mux2_1
XANTENNA_38 _11634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_49 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05382_ _10465_/Q _10464_/Q _05382_/S vssd1 vssd1 vccd1 vccd1 _05384_/C sky130_fd_sc_hd__mux2_1
XFILLER_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07121_ _10318_/Q _07126_/B _07186_/S _07314_/B vssd1 vssd1 vccd1 vccd1 _10318_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07052_ _07052_/A _10028_/A vssd1 vssd1 vccd1 vccd1 _07052_/X sky130_fd_sc_hd__and2_4
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06003_ _10938_/Q _10061_/A _06630_/B1 _11014_/Q vssd1 vssd1 vccd1 vccd1 _06003_/X
+ sky130_fd_sc_hd__o22a_1
Xoutput123 _05680_/X vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_4
Xoutput134 _11614_/Q vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_4
Xoutput145 _10213_/Q vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__buf_4
Xoutput156 _10221_/Q vssd1 vssd1 vccd1 vccd1 ram_val_out[3] sky130_fd_sc_hd__buf_4
XFILLER_138_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput167 _09959_/A vssd1 vssd1 vccd1 vccd1 rom_csb sky130_fd_sc_hd__buf_4
XFILLER_82_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput178 _06892_/A vssd1 vssd1 vccd1 vccd1 wb_rom_web sky130_fd_sc_hd__buf_4
XFILLER_141_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput189 _05495_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_4
XFILLER_138_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07954_ _07013_/X _10796_/Q _07961_/S vssd1 vssd1 vccd1 vccd1 _10796_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06905_ _10088_/A1 _06903_/X _06904_/X _06990_/C1 vssd1 vssd1 vccd1 vccd1 _10193_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07885_ _10761_/Q _07901_/B vssd1 vssd1 vccd1 vccd1 _07885_/X sky130_fd_sc_hd__or2_1
XFILLER_96_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09624_ _10801_/Q _09571_/A _09950_/B1 _10722_/Q vssd1 vssd1 vccd1 vccd1 _09626_/C
+ sky130_fd_sc_hd__a22o_1
X_06836_ _11474_/Q _07153_/A _06835_/X _06878_/C1 vssd1 vssd1 vccd1 vccd1 _06836_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09555_ _05074_/Y _09692_/B _09673_/B _09554_/Y _09959_/A vssd1 vssd1 vccd1 vccd1
+ _11629_/D sky130_fd_sc_hd__a221oi_1
Xclkbuf_leaf_37_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11735_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_06767_ _06762_/X _06763_/X _06766_/X _06761_/X vssd1 vssd1 vccd1 vccd1 _06767_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_52_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08506_ _09082_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08506_/X sky130_fd_sc_hd__or2_4
X_05718_ _10963_/Q _05549_/Y _05603_/Y _10959_/Q vssd1 vssd1 vccd1 vccd1 _05727_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_145_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09486_ _09522_/B _09515_/B _09515_/C vssd1 vssd1 vccd1 vccd1 _09486_/X sky130_fd_sc_hd__or3_1
XFILLER_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06698_ _11330_/Q _06738_/A2 _06739_/A2 _11302_/Q _06718_/C1 vssd1 vssd1 vccd1 vccd1
+ _06698_/X sky130_fd_sc_hd__o221a_1
XFILLER_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08437_ _08437_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08437_/Y sky130_fd_sc_hd__nand2_2
XFILLER_145_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05649_ _11291_/Q _05537_/Y _05573_/Y _11294_/Q _05648_/X vssd1 vssd1 vccd1 vccd1
+ _05655_/C sky130_fd_sc_hd__a221o_1
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08368_ _09256_/A1 _11026_/Q _08439_/B vssd1 vssd1 vccd1 vccd1 _08369_/B sky130_fd_sc_hd__mux2_1
XFILLER_149_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07319_ _10426_/Q _07302_/Y _07305_/Y _07318_/X vssd1 vssd1 vccd1 vccd1 _10426_/D
+ sky130_fd_sc_hd__o22a_1
X_08299_ _09248_/A _08471_/B _09037_/C vssd1 vssd1 vccd1 vccd1 _08840_/B sky130_fd_sc_hd__and3_4
X_10330_ _11710_/CLK _10330_/D vssd1 vssd1 vccd1 vccd1 _10330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10261_ _11808_/CLK _10261_/D vssd1 vssd1 vccd1 vccd1 _10261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10192_ _09497_/A _09486_/X _09528_/B _10191_/X _09825_/A vssd1 vssd1 vccd1 vccd1
+ _11812_/D sky130_fd_sc_hd__o311a_1
XFILLER_152_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout350 _07643_/C vssd1 vssd1 vccd1 vccd1 _08560_/C sky130_fd_sc_hd__buf_4
Xfanout361 _10180_/B vssd1 vssd1 vccd1 vccd1 _10108_/B sky130_fd_sc_hd__buf_4
Xfanout372 _09206_/A vssd1 vssd1 vccd1 vccd1 _09227_/A sky130_fd_sc_hd__buf_6
XFILLER_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout383 _08439_/A vssd1 vssd1 vccd1 vccd1 _08427_/A sky130_fd_sc_hd__buf_6
XFILLER_98_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout394 _09228_/A vssd1 vssd1 vccd1 vccd1 _09192_/A sky130_fd_sc_hd__buf_6
XFILLER_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _11719_/CLK _11715_/D vssd1 vssd1 vccd1 vccd1 _11715_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11646_ _11665_/CLK _11646_/D vssd1 vssd1 vccd1 vccd1 _11646_/Q sky130_fd_sc_hd__dfxtp_1
Xinput14 rom_value[13] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
Xinput25 rom_value[23] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_2
Xinput36 rom_value[4] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_2
X_11577_ _11650_/CLK _11577_/D vssd1 vssd1 vccd1 vccd1 _11577_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 wb_rom_val[14] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_2
XFILLER_7_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput58 wb_rom_val[24] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_4
X_10528_ _11720_/CLK _10528_/D vssd1 vssd1 vccd1 vccd1 _10528_/Q sky130_fd_sc_hd__dfxtp_1
Xinput69 wb_rom_val[5] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_2
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10459_ _11308_/CLK _10459_/D vssd1 vssd1 vccd1 vccd1 _10459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07670_ _10631_/Q _07665_/S _07249_/S _07040_/B vssd1 vssd1 vccd1 vccd1 _10631_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_93_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06621_ _06535_/A _06620_/X _06619_/X _06664_/C1 vssd1 vssd1 vccd1 vccd1 _06621_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09340_ _11524_/Q _09326_/X _09339_/X vssd1 vssd1 vccd1 vccd1 _11524_/D sky130_fd_sc_hd__a21o_1
X_06552_ _06552_/A _06552_/B _06552_/C vssd1 vssd1 vccd1 vccd1 _06552_/X sky130_fd_sc_hd__and3_1
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05503_ _10248_/Q input60/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05503_/X sky130_fd_sc_hd__mux2_2
X_09271_ _09271_/A _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09271_/X sky130_fd_sc_hd__or3_4
XFILLER_61_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06483_ _10485_/Q _08649_/A _06481_/X _06482_/X vssd1 vssd1 vccd1 vccd1 _06483_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_61_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08222_ _08839_/A _08222_/B vssd1 vssd1 vccd1 vccd1 _10945_/D sky130_fd_sc_hd__or2_1
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05434_ _05434_/A _05434_/B vssd1 vssd1 vccd1 vccd1 _05434_/Y sky130_fd_sc_hd__nor2_8
XFILLER_147_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08153_ _09985_/A1 _08162_/S _08152_/X _07011_/B vssd1 vssd1 vccd1 vccd1 _10902_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05365_ _11278_/Q _11277_/Q _09680_/B vssd1 vssd1 vccd1 vccd1 _05367_/C sky130_fd_sc_hd__mux2_1
XFILLER_147_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07104_ _07104_/A _10028_/A vssd1 vssd1 vccd1 vccd1 _07333_/B sky130_fd_sc_hd__and2_4
X_08084_ _08761_/A _08084_/B vssd1 vssd1 vccd1 vccd1 _10867_/D sky130_fd_sc_hd__or2_1
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05296_ _05296_/A _05296_/B _05296_/C _05296_/D vssd1 vssd1 vccd1 vccd1 _05302_/A
+ sky130_fd_sc_hd__or4_4
X_07035_ _10276_/Q _07000_/Y _07034_/X _07000_/B _07333_/A vssd1 vssd1 vccd1 vccd1
+ _10276_/D sky130_fd_sc_hd__a221o_1
XFILLER_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08986_ _09285_/A1 _08972_/X _08985_/X _09279_/C1 vssd1 vssd1 vccd1 vccd1 _11345_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07937_ _07143_/A _10786_/Q _09221_/C vssd1 vssd1 vccd1 vccd1 _07938_/B sky130_fd_sc_hd__mux2_1
XFILLER_112_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07868_ _09214_/A _07871_/S _07867_/X _07868_/C1 vssd1 vssd1 vccd1 vccd1 _10752_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06819_ _10333_/Q _06856_/A2 _06685_/B _11720_/Q vssd1 vssd1 vccd1 vccd1 _06819_/X
+ sky130_fd_sc_hd__o22a_1
X_09607_ _10632_/Q _09572_/A _09571_/D _10621_/Q _09606_/X vssd1 vssd1 vccd1 vccd1
+ _09617_/B sky130_fd_sc_hd__a221o_1
X_07799_ _08883_/A1 _10707_/Q _09200_/S vssd1 vssd1 vccd1 vccd1 _07800_/B sky130_fd_sc_hd__mux2_1
XFILLER_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09538_ _09538_/A _09538_/B _09538_/C _09538_/D vssd1 vssd1 vccd1 vccd1 _09538_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_19_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09469_ input38/X _09442_/X _09468_/X vssd1 vssd1 vccd1 vccd1 _09470_/B sky130_fd_sc_hd__o21ai_1
XFILLER_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11500_ _11800_/CLK _11500_/D vssd1 vssd1 vccd1 vccd1 _11500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11431_ _11431_/CLK _11431_/D vssd1 vssd1 vccd1 vccd1 _11431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11362_ _11366_/CLK _11362_/D vssd1 vssd1 vccd1 vccd1 _11362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10313_ _10812_/CLK _10313_/D vssd1 vssd1 vccd1 vccd1 _10313_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11293_ _11325_/CLK _11293_/D vssd1 vssd1 vccd1 vccd1 _11293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10244_ _11712_/CLK _10244_/D vssd1 vssd1 vccd1 vccd1 _10244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10175_ _10175_/A1 _10159_/X _10174_/X _10175_/C1 vssd1 vssd1 vccd1 vccd1 _11799_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11629_ _11629_/CLK _11629_/D vssd1 vssd1 vccd1 vccd1 _11629_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05150_ _10940_/Q _10939_/Q _05372_/S vssd1 vssd1 vccd1 vccd1 _05151_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05081_ _09680_/B vssd1 vssd1 vccd1 vccd1 _06941_/A sky130_fd_sc_hd__inv_2
XFILLER_100_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _11278_/Q _08840_/B vssd1 vssd1 vccd1 vccd1 _08840_/X sky130_fd_sc_hd__or2_1
XFILLER_135_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08771_ _08771_/A _08771_/B vssd1 vssd1 vccd1 vccd1 _11241_/D sky130_fd_sc_hd__or2_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05983_ _10684_/Q _07203_/A _05979_/X _05982_/X vssd1 vssd1 vccd1 vccd1 _05983_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_85_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07722_ _10662_/Q _07750_/B vssd1 vssd1 vccd1 vccd1 _07722_/X sky130_fd_sc_hd__or2_1
XFILLER_38_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07653_ _08441_/B2 _10617_/Q _07655_/S vssd1 vssd1 vccd1 vccd1 _10617_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06604_ _10708_/Q _09059_/A _09109_/A _10543_/Q _06603_/X vssd1 vssd1 vccd1 vccd1
+ _06604_/X sky130_fd_sc_hd__a221o_1
XFILLER_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07584_ _07812_/A _07584_/B vssd1 vssd1 vccd1 vccd1 _10575_/D sky130_fd_sc_hd__or2_1
XFILLER_0_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09323_ _09323_/A0 _11516_/Q _09324_/S vssd1 vssd1 vccd1 vccd1 _11516_/D sky130_fd_sc_hd__mux2_1
X_06535_ _06535_/A _06535_/B vssd1 vssd1 vccd1 vccd1 _06535_/X sky130_fd_sc_hd__or2_1
XFILLER_90_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ _11480_/Q _09266_/B vssd1 vssd1 vccd1 vccd1 _09254_/X sky130_fd_sc_hd__or2_1
XFILLER_139_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06466_ _10606_/Q _06635_/B1 _10119_/A _11777_/Q _06465_/X vssd1 vssd1 vccd1 vccd1
+ _06467_/C sky130_fd_sc_hd__o221a_1
XFILLER_107_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08205_ _10937_/Q _08902_/C vssd1 vssd1 vccd1 vccd1 _08205_/X sky130_fd_sc_hd__or2_1
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05417_ _05417_/A _05417_/B _05417_/C _05417_/D vssd1 vssd1 vccd1 vccd1 _05423_/A
+ sky130_fd_sc_hd__or4_4
X_09185_ _07812_/A _09184_/X _09227_/A vssd1 vssd1 vccd1 vccd1 _11437_/D sky130_fd_sc_hd__o21a_1
X_06397_ _10469_/Q _06642_/A2 _06393_/X _06396_/X vssd1 vssd1 vccd1 vccd1 _06397_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08136_ _10894_/Q _08637_/C vssd1 vssd1 vccd1 vccd1 _08136_/X sky130_fd_sc_hd__or2_1
X_05348_ _11138_/Q _11137_/Q _05392_/S vssd1 vssd1 vccd1 vccd1 _05354_/B sky130_fd_sc_hd__mux2_1
XFILLER_88_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08067_ _08838_/A0 _10859_/Q _08427_/B vssd1 vssd1 vccd1 vccd1 _08068_/B sky130_fd_sc_hd__mux2_1
X_05279_ _10817_/Q _10816_/Q _05394_/S vssd1 vssd1 vccd1 vccd1 _05280_/D sky130_fd_sc_hd__mux2_1
XFILLER_150_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07018_ _07018_/A _07018_/B vssd1 vssd1 vccd1 vccd1 _07018_/X sky130_fd_sc_hd__and2_1
XFILLER_134_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_52_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11067_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08969_ _11337_/Q _08969_/A1 _08970_/S vssd1 vssd1 vccd1 vccd1 _11337_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10931_ _11584_/CLK _10931_/D vssd1 vssd1 vccd1 vccd1 _10931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10862_ _11628_/CLK _10862_/D vssd1 vssd1 vccd1 vccd1 _10862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _11005_/CLK _10793_/D vssd1 vssd1 vccd1 vccd1 _10793_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11414_ _11792_/CLK _11414_/D vssd1 vssd1 vccd1 vccd1 _11414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11345_ _11495_/CLK _11345_/D vssd1 vssd1 vccd1 vccd1 _11345_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11276_ _11604_/CLK _11276_/D vssd1 vssd1 vccd1 vccd1 _11276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10227_ _11233_/CLK _10227_/D vssd1 vssd1 vccd1 vccd1 _10227_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10158_ _10158_/A _10158_/B _10158_/C vssd1 vssd1 vccd1 vccd1 _10176_/B sky130_fd_sc_hd__and3_4
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10089_ _11746_/Q _10087_/X _10088_/X vssd1 vssd1 vccd1 vccd1 _11746_/D sky130_fd_sc_hd__a21o_1
XFILLER_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06320_ _10791_/Q _06540_/A2 _06540_/B1 _10905_/Q vssd1 vssd1 vccd1 vccd1 _06320_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06251_ _11184_/Q _06470_/A2 _06639_/B1 _10815_/Q vssd1 vssd1 vccd1 vccd1 _06255_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_50_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05202_ _05419_/S _11067_/Q _11066_/Q _09679_/B _05196_/X vssd1 vssd1 vccd1 vccd1
+ _05204_/C sky130_fd_sc_hd__a221oi_2
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06182_ _11762_/Q _10108_/A _06180_/X _06181_/X vssd1 vssd1 vccd1 vccd1 _06182_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05133_ _10930_/Q _10929_/Q _05394_/S vssd1 vssd1 vccd1 vccd1 _05134_/D sky130_fd_sc_hd__mux2_1
X_09941_ _10684_/Q _09566_/C _09572_/C _10374_/Q vssd1 vssd1 vccd1 vccd1 _09941_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout905 _05095_/Y vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__buf_12
Xfanout916 _07689_/B vssd1 vssd1 vccd1 vccd1 _06265_/C1 sky130_fd_sc_hd__buf_6
Xfanout927 _09393_/A0 vssd1 vssd1 vccd1 vccd1 _10110_/A0 sky130_fd_sc_hd__clkbuf_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _10577_/Q _09872_/A2 _09872_/B1 _10559_/Q vssd1 vssd1 vccd1 vccd1 _09872_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 _08893_/A1 vssd1 vssd1 vccd1 vccd1 _07031_/A sky130_fd_sc_hd__buf_6
XFILLER_135_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout949 _08939_/A1 vssd1 vssd1 vccd1 vccd1 _08853_/A1 sky130_fd_sc_hd__buf_6
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08833_/A _08823_/B vssd1 vssd1 vccd1 vccd1 _11269_/D sky130_fd_sc_hd__or2_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_7__f_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_7__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _09256_/A1 _11234_/Q _08760_/S vssd1 vssd1 vccd1 vccd1 _08755_/B sky130_fd_sc_hd__mux2_1
XFILLER_100_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05966_ _11759_/Q _10108_/A _05964_/X _05965_/X vssd1 vssd1 vccd1 vccd1 _05966_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07705_ _10653_/Q _07694_/Y _07696_/Y _07318_/X vssd1 vssd1 vccd1 vccd1 _10653_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _09172_/A1 _11197_/Q _08695_/S vssd1 vssd1 vccd1 vccd1 _08686_/B sky130_fd_sc_hd__mux2_1
X_05897_ _11668_/Q _09965_/A _06284_/B1 _10993_/Q vssd1 vssd1 vccd1 vccd1 _05897_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07636_ _10605_/Q _07100_/X _07637_/S vssd1 vssd1 vccd1 vccd1 _10605_/D sky130_fd_sc_hd__mux2_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07567_ _08883_/A1 _10567_/Q _07589_/S vssd1 vssd1 vccd1 vccd1 _07568_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09306_ _10172_/A1 _09310_/B _10178_/B1 vssd1 vssd1 vccd1 vccd1 _09306_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06518_ _10776_/Q _06646_/A2 _08971_/A _10566_/Q vssd1 vssd1 vccd1 vccd1 _06518_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07498_ _10013_/A0 _07513_/S _07497_/X _07868_/C1 vssd1 vssd1 vccd1 vccd1 _10533_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09237_ _09237_/A0 _11470_/Q _09240_/S vssd1 vssd1 vccd1 vccd1 _09237_/X sky130_fd_sc_hd__mux2_1
X_06449_ _07081_/A _06420_/X _06431_/X _06448_/X vssd1 vssd1 vccd1 vccd1 _06449_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09168_ _10172_/A1 _09154_/X _09167_/X _09168_/C1 vssd1 vssd1 vccd1 vccd1 _11428_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08119_ _08193_/A _08119_/B vssd1 vssd1 vccd1 vccd1 _10886_/D sky130_fd_sc_hd__or2_1
X_09099_ _11397_/Q _09099_/B vssd1 vssd1 vccd1 vccd1 _09099_/X sky130_fd_sc_hd__or2_1
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11130_ _11777_/CLK _11130_/D vssd1 vssd1 vccd1 vccd1 _11130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11061_ _11067_/CLK _11061_/D vssd1 vssd1 vccd1 vccd1 _11061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10012_ _10026_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _11696_/D sky130_fd_sc_hd__or2_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10914_ _11780_/CLK _10914_/D vssd1 vssd1 vccd1 vccd1 _10914_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10845_ _11308_/CLK _10845_/D vssd1 vssd1 vccd1 vccd1 _10845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10776_ _11450_/CLK _10776_/D vssd1 vssd1 vccd1 vccd1 _10776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ _11330_/CLK _11328_/D vssd1 vssd1 vccd1 vccd1 _11328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11259_ _11770_/CLK _11259_/D vssd1 vssd1 vccd1 vccd1 _11259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05820_ _06892_/A _05820_/B vssd1 vssd1 vccd1 vccd1 _06883_/B sky130_fd_sc_hd__nand2_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05751_ _05751_/A _05751_/B _11867_/A vssd1 vssd1 vccd1 vccd1 _05751_/X sky130_fd_sc_hd__or3b_4
XFILLER_35_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08470_ _11086_/Q _08467_/S _08469_/X _08578_/A vssd1 vssd1 vccd1 vccd1 _11086_/D
+ sky130_fd_sc_hd__o211a_1
X_05682_ _11154_/Q _05531_/Y _05591_/Y _11170_/Q _05681_/X vssd1 vssd1 vccd1 vccd1
+ _05692_/A sky130_fd_sc_hd__a221o_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07421_ _07025_/A _10487_/Q _07437_/S vssd1 vssd1 vccd1 vccd1 _07422_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07352_ _07939_/A _08560_/C _07847_/C vssd1 vssd1 vccd1 vccd1 _07353_/B sky130_fd_sc_hd__and3_4
XFILLER_17_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06303_ _11466_/Q _07152_/A _06805_/B1 _10499_/Q _06302_/X vssd1 vssd1 vccd1 vccd1
+ _06303_/X sky130_fd_sc_hd__o221a_1
XFILLER_17_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07283_ _08423_/A1 _10410_/Q _09184_/S vssd1 vssd1 vccd1 vccd1 _07284_/B sky130_fd_sc_hd__mux2_1
X_09022_ _10183_/A0 _09016_/X _09021_/X _09022_/C1 vssd1 vssd1 vccd1 vccd1 _11361_/D
+ sky130_fd_sc_hd__o211a_1
X_06234_ _11870_/A _06223_/X _06232_/X _06233_/X _08243_/A vssd1 vssd1 vccd1 vccd1
+ _06234_/X sky130_fd_sc_hd__o221a_2
XFILLER_148_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06165_ _10421_/Q _06541_/A2 _06540_/A2 _10790_/Q _06164_/X vssd1 vssd1 vccd1 vccd1
+ _06165_/X sky130_fd_sc_hd__o221a_1
XFILLER_105_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05116_ _11176_/Q _10301_/Q _05396_/S vssd1 vssd1 vccd1 vccd1 _05118_/C sky130_fd_sc_hd__mux2_1
XFILLER_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06096_ _11691_/Q _09998_/A _06924_/A _11738_/Q _06344_/C1 vssd1 vssd1 vccd1 vccd1
+ _06096_/X sky130_fd_sc_hd__o221a_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09924_ _10361_/Q _09566_/D _09573_/D _10480_/Q _09923_/X vssd1 vssd1 vccd1 vccd1
+ _09925_/D sky130_fd_sc_hd__a221o_1
Xfanout702 _05418_/S vssd1 vssd1 vccd1 vccd1 _09539_/B sky130_fd_sc_hd__buf_8
XFILLER_104_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout713 _05786_/Y vssd1 vssd1 vccd1 vccd1 _07081_/A sky130_fd_sc_hd__buf_6
Xfanout724 _06540_/B1 vssd1 vssd1 vccd1 vccd1 _06903_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_63_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout735 _08765_/A vssd1 vssd1 vccd1 vccd1 _09110_/A sky130_fd_sc_hd__clkbuf_8
Xfanout746 fanout755/X vssd1 vssd1 vccd1 vccd1 _10010_/A sky130_fd_sc_hd__buf_4
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout757 _06674_/A2 vssd1 vssd1 vccd1 vccd1 _06857_/B1 sky130_fd_sc_hd__buf_6
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _10697_/Q _09874_/A2 _09567_/C _10704_/Q vssd1 vssd1 vccd1 vccd1 _09855_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout768 _05748_/Y vssd1 vssd1 vccd1 vccd1 _10136_/A sky130_fd_sc_hd__buf_12
XFILLER_100_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout779 _06538_/B1 vssd1 vssd1 vccd1 vccd1 _06453_/B1 sky130_fd_sc_hd__buf_4
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _11259_/Q _07092_/A _08820_/S vssd1 vssd1 vccd1 vccd1 _08807_/B sky130_fd_sc_hd__mux2_1
XFILLER_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06998_ _06998_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _07000_/B sky130_fd_sc_hd__nor2_8
XFILLER_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09786_ _11649_/Q _08950_/B _09785_/X _09407_/A vssd1 vssd1 vccd1 vccd1 _11649_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ _08749_/A _08737_/B vssd1 vssd1 vccd1 vccd1 _11225_/D sky130_fd_sc_hd__or2_1
X_05949_ _05668_/X _06622_/A2 _05886_/X _06886_/A2 vssd1 vssd1 vccd1 vccd1 _05950_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 _09292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _06194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_128 _09214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _05179_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _08668_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08683_/S sky130_fd_sc_hd__or2_4
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ _10594_/Q _07613_/Y _07614_/Y _07016_/X vssd1 vssd1 vccd1 vccd1 _10594_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _09364_/A1 _11154_/Q _08621_/S vssd1 vssd1 vccd1 vccd1 _08600_/B sky130_fd_sc_hd__mux2_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10630_ _11745_/CLK _10630_/D vssd1 vssd1 vccd1 vccd1 _10630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10561_ _11622_/CLK _10561_/D vssd1 vssd1 vccd1 vccd1 _10561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10492_ _11719_/CLK _10492_/D vssd1 vssd1 vccd1 vccd1 _10492_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11113_ _11572_/CLK _11113_/D vssd1 vssd1 vccd1 vccd1 _11113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11044_ _11683_/CLK _11044_/D vssd1 vssd1 vccd1 vccd1 _11044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10828_ _11634_/CLK _10828_/D vssd1 vssd1 vccd1 vccd1 _10828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10759_ _11470_/CLK _10759_/D vssd1 vssd1 vccd1 vccd1 _10759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07970_ input103/X _10808_/Q _07970_/S vssd1 vssd1 vccd1 vccd1 _07970_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06921_ _10201_/Q _06903_/X _06920_/X vssd1 vssd1 vccd1 vccd1 _10201_/D sky130_fd_sc_hd__a21o_1
XFILLER_45_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06852_ _06852_/A1 _10249_/Q _06852_/A3 _06743_/X _06851_/X vssd1 vssd1 vccd1 vccd1
+ _06852_/X sky130_fd_sc_hd__a32o_1
XFILLER_45_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09640_ _09820_/A _09640_/B _09640_/C vssd1 vssd1 vccd1 vccd1 _09640_/X sky130_fd_sc_hd__and3b_1
Xclkbuf_leaf_109_wb_clk_i clkbuf_4_10__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10548_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05803_ _11135_/Q _10010_/A _05799_/X _05802_/X vssd1 vssd1 vccd1 vccd1 _05803_/X
+ sky130_fd_sc_hd__o211a_1
X_09571_ _09571_/A _09571_/B _09571_/C _09571_/D vssd1 vssd1 vccd1 vccd1 _09574_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06783_ _06853_/A1 _10244_/Q _06853_/A3 _06782_/X _05730_/Y vssd1 vssd1 vccd1 vccd1
+ _06783_/X sky130_fd_sc_hd__a32o_1
XFILLER_36_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08522_ _08987_/A1 _08537_/S _08521_/X _08937_/C1 vssd1 vssd1 vccd1 vccd1 _11110_/D
+ sky130_fd_sc_hd__o211a_1
X_05734_ _05819_/A _06892_/B vssd1 vssd1 vccd1 vccd1 _05734_/X sky130_fd_sc_hd__or2_4
XFILLER_36_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08453_ _11074_/Q _08459_/S _07626_/S _07617_/B vssd1 vssd1 vccd1 vccd1 _11074_/D
+ sky130_fd_sc_hd__o22a_1
X_05665_ _11254_/Q _05561_/Y _05585_/Y _11253_/Q _05664_/X vssd1 vssd1 vccd1 vccd1
+ _05668_/C sky130_fd_sc_hd__a221o_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07404_ _10020_/A _07404_/B vssd1 vssd1 vccd1 vccd1 _10478_/D sky130_fd_sc_hd__or2_1
XFILLER_17_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08384_ _08669_/A0 _11033_/Q _08404_/S vssd1 vssd1 vccd1 vccd1 _08385_/B sky130_fd_sc_hd__mux2_1
X_05596_ _05626_/A2 _11484_/Q _11479_/Q _05630_/B1 _05595_/X vssd1 vssd1 vccd1 vccd1
+ _05597_/B sky130_fd_sc_hd__a221o_4
XFILLER_108_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07335_ _08322_/A _07335_/B vssd1 vssd1 vccd1 vccd1 _07335_/X sky130_fd_sc_hd__or2_4
XFILLER_91_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07266_ _07920_/A _07266_/B vssd1 vssd1 vccd1 vccd1 _10401_/D sky130_fd_sc_hd__or2_1
X_09005_ _11354_/Q _09013_/B vssd1 vssd1 vccd1 vccd1 _09005_/X sky130_fd_sc_hd__or2_1
X_06217_ _11683_/Q _08594_/A _06213_/X _06216_/X vssd1 vssd1 vccd1 vccd1 _06217_/X
+ sky130_fd_sc_hd__o211a_1
X_07197_ _07070_/A _07191_/B _07192_/A _10359_/Q _07333_/A vssd1 vssd1 vccd1 vccd1
+ _10359_/D sky130_fd_sc_hd__a221o_1
XFILLER_133_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06148_ _10879_/Q _06513_/A2 _06636_/A2 _10927_/Q _07083_/B vssd1 vssd1 vccd1 vccd1
+ _06151_/B sky130_fd_sc_hd__o221a_1
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06079_ _05816_/A _06017_/Y _05820_/B vssd1 vssd1 vccd1 vccd1 _06079_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_120_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout510 _06899_/X vssd1 vssd1 vccd1 vccd1 fanout510/X sky130_fd_sc_hd__buf_8
XFILLER_120_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout521 _07664_/A vssd1 vssd1 vccd1 vccd1 _07420_/A sky130_fd_sc_hd__clkbuf_4
Xfanout532 _10150_/B1 vssd1 vssd1 vccd1 vccd1 _10156_/B1 sky130_fd_sc_hd__buf_4
X_09907_ _09907_/A _09907_/B _09907_/C _09907_/D vssd1 vssd1 vccd1 vccd1 _09908_/B
+ sky130_fd_sc_hd__or4_4
Xfanout543 fanout555/X vssd1 vssd1 vccd1 vccd1 _10020_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout554 fanout555/X vssd1 vssd1 vccd1 vccd1 _07790_/A sky130_fd_sc_hd__buf_4
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout565 _08773_/A vssd1 vssd1 vccd1 vccd1 fanout565/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout576 fanout578/X vssd1 vssd1 vccd1 vccd1 _08869_/A sky130_fd_sc_hd__buf_4
XFILLER_47_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ _11457_/Q _09881_/A2 _09878_/A2 _11458_/Q vssd1 vssd1 vccd1 vccd1 _09838_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout587 _05734_/X vssd1 vssd1 vccd1 vccd1 _06576_/A sky130_fd_sc_hd__buf_4
XFILLER_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout598 _09015_/B vssd1 vssd1 vccd1 vccd1 _08649_/B sky130_fd_sc_hd__buf_6
XFILLER_111_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09769_ input9/X _09740_/Y _09768_/X vssd1 vssd1 vccd1 vccd1 _09769_/X sky130_fd_sc_hd__a21o_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _11800_/CLK _11800_/D vssd1 vssd1 vccd1 vccd1 _11800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11765_/CLK _11731_/D vssd1 vssd1 vccd1 vccd1 _11731_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11663_/CLK _11662_/D vssd1 vssd1 vccd1 vccd1 _11662_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10613_ _10932_/CLK _10613_/D vssd1 vssd1 vccd1 vccd1 _10613_/Q sky130_fd_sc_hd__dfxtp_1
X_11593_ _11652_/CLK _11593_/D vssd1 vssd1 vccd1 vccd1 _11593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10544_ _10548_/CLK _10544_/D vssd1 vssd1 vccd1 vccd1 _10544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10475_ _10725_/CLK _10475_/D vssd1 vssd1 vccd1 vccd1 _10475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11641_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11027_ _11067_/CLK _11027_/D vssd1 vssd1 vccd1 vccd1 _11027_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05450_ _10676_/Q _09572_/B _09573_/C _10674_/Q _05437_/X vssd1 vssd1 vccd1 vccd1
+ _05451_/D sky130_fd_sc_hd__a221o_1
XFILLER_92_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _06205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _07008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 _11718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05381_ _10467_/Q _10466_/Q _05414_/S vssd1 vssd1 vccd1 vccd1 _05384_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07120_ _10317_/Q _07135_/A2 _07123_/B1 _07022_/B vssd1 vssd1 vccd1 vccd1 _10317_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07051_ _10282_/Q _07047_/B _07490_/S _07227_/B vssd1 vssd1 vccd1 vccd1 _10282_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_51_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06002_ _11056_/Q _08054_/A _08123_/A _10890_/Q _06392_/C1 vssd1 vssd1 vccd1 vccd1
+ _06002_/X sky130_fd_sc_hd__o221a_1
XFILLER_127_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput124 _05692_/X vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_4
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput135 _11615_/Q vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_4
Xoutput146 _11569_/Q vssd1 vssd1 vccd1 vccd1 ram_addr[0] sky130_fd_sc_hd__buf_4
Xoutput157 _05475_/X vssd1 vssd1 vccd1 vccd1 ram_we sky130_fd_sc_hd__buf_4
Xoutput168 _11866_/X vssd1 vssd1 vccd1 vccd1 wb_rom_adrb[0] sky130_fd_sc_hd__buf_4
Xoutput179 _10254_/Q vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_4
XFILLER_47_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07953_ _08326_/B2 _10795_/Q _07956_/S vssd1 vssd1 vccd1 vccd1 _10795_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06904_ _10193_/Q _06922_/B vssd1 vssd1 vccd1 vccd1 _06904_/X sky130_fd_sc_hd__or2_1
X_07884_ _08893_/A1 _07970_/S _07883_/X _07884_/C1 vssd1 vssd1 vccd1 vccd1 _10760_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09623_ _10724_/Q _09947_/A2 _09568_/D _10795_/Q vssd1 vssd1 vccd1 vccd1 _09626_/B
+ sky130_fd_sc_hd__a22o_1
X_06835_ _11460_/Q _06875_/A2 _06877_/B1 _10580_/Q _06834_/X vssd1 vssd1 vccd1 vccd1
+ _06835_/X sky130_fd_sc_hd__o221a_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06766_ _10351_/Q _06766_/A2 _06765_/X _06878_/C1 vssd1 vssd1 vccd1 vccd1 _06766_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09554_ _09554_/A _09554_/B vssd1 vssd1 vccd1 vccd1 _09554_/Y sky130_fd_sc_hd__nor2_4
XFILLER_110_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05717_ _10972_/Q _05543_/Y _05615_/Y _10968_/Q vssd1 vssd1 vccd1 vccd1 _05727_/A
+ sky130_fd_sc_hd__a22o_1
X_08505_ _09082_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08545_/B sky130_fd_sc_hd__nor2_8
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09485_ _09522_/B _09504_/B vssd1 vssd1 vccd1 vccd1 _09485_/X sky130_fd_sc_hd__and2b_1
X_06697_ _11120_/Q _06737_/A2 _06697_/B1 _11256_/Q vssd1 vssd1 vccd1 vccd1 _06697_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_93_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08436_ _08902_/B _08438_/B vssd1 vssd1 vccd1 vccd1 _08436_/Y sky130_fd_sc_hd__nor2_2
X_05648_ _11304_/Q _05518_/Y _05524_/Y _11295_/Q vssd1 vssd1 vccd1 vccd1 _05648_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_77_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11325_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08367_ _10142_/A1 _08439_/B _08366_/X _08662_/C1 vssd1 vssd1 vccd1 vccd1 _11025_/D
+ sky130_fd_sc_hd__o211a_1
X_05579_ _05579_/A _05579_/B vssd1 vssd1 vccd1 vccd1 _05579_/Y sky130_fd_sc_hd__nor2_8
XFILLER_149_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07318_ _07318_/A _07318_/B vssd1 vssd1 vccd1 vccd1 _07318_/X sky130_fd_sc_hd__or2_4
X_08298_ _10984_/Q _08901_/A1 _08298_/S vssd1 vssd1 vccd1 vccd1 _10984_/D sky130_fd_sc_hd__mux2_1
X_07249_ _07248_/X _10393_/Q _07249_/S vssd1 vssd1 vccd1 vccd1 _10393_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ _11755_/CLK _10260_/D vssd1 vssd1 vccd1 vccd1 _10260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10191_ _09525_/A _09485_/X _09489_/C _11812_/Q vssd1 vssd1 vccd1 vccd1 _10191_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout340 _08951_/X vssd1 vssd1 vccd1 vccd1 _09959_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout351 _08471_/B vssd1 vssd1 vccd1 vccd1 _08649_/C sky130_fd_sc_hd__buf_6
Xfanout362 _09407_/B vssd1 vssd1 vccd1 vccd1 _09475_/A sky130_fd_sc_hd__clkbuf_4
Xfanout373 _07012_/Y vssd1 vssd1 vccd1 vccd1 _09206_/A sky130_fd_sc_hd__buf_12
XFILLER_115_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout384 _07004_/Y vssd1 vssd1 vccd1 vccd1 _08439_/A sky130_fd_sc_hd__buf_12
XFILLER_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout395 _07599_/A vssd1 vssd1 vccd1 vccd1 _09228_/A sky130_fd_sc_hd__buf_6
XFILLER_115_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11720_/CLK _11714_/D vssd1 vssd1 vccd1 vccd1 _11714_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _11665_/CLK _11645_/D vssd1 vssd1 vccd1 vccd1 _11645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 rom_value[14] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
Xinput26 rom_value[24] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_2
X_11576_ _11650_/CLK _11576_/D vssd1 vssd1 vccd1 vccd1 _11576_/Q sky130_fd_sc_hd__dfxtp_4
Xinput37 rom_value[5] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_2
Xinput48 wb_rom_val[15] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_2
XFILLER_156_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput59 wb_rom_val[25] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10527_ _11711_/CLK _10527_/D vssd1 vssd1 vccd1 vccd1 _10527_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10458_ _11308_/CLK _10458_/D vssd1 vssd1 vccd1 vccd1 _10458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10389_ _11477_/CLK _10389_/D vssd1 vssd1 vccd1 vccd1 _10389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06620_ _06663_/A _10236_/Q vssd1 vssd1 vccd1 vccd1 _06620_/X sky130_fd_sc_hd__and2_1
XFILLER_53_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06551_ _11266_/Q _06635_/B1 _10119_/A _11779_/Q _06550_/X vssd1 vssd1 vccd1 vccd1
+ _06552_/C sky130_fd_sc_hd__o221a_1
XFILLER_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05502_ _10247_/Q input59/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05502_/X sky130_fd_sc_hd__mux2_1
X_09270_ _10086_/A _09270_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09288_/B sky130_fd_sc_hd__and3_4
X_06482_ _10625_/Q _07939_/A _08286_/A _10724_/Q vssd1 vssd1 vccd1 vccd1 _06482_/X
+ sky130_fd_sc_hd__a22o_1
X_08221_ _08834_/A0 _10945_/Q _08225_/S vssd1 vssd1 vccd1 vccd1 _08222_/B sky130_fd_sc_hd__mux2_1
X_05433_ _05433_/A _05433_/B _05433_/C _05433_/D vssd1 vssd1 vccd1 vccd1 _05434_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _10902_/Q _08164_/B vssd1 vssd1 vccd1 vccd1 _08152_/X sky130_fd_sc_hd__or2_1
X_05364_ _11276_/Q _11275_/Q _09680_/C vssd1 vssd1 vccd1 vccd1 _05367_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07103_ _10307_/Q _08901_/A1 _07109_/S vssd1 vssd1 vccd1 vccd1 _10307_/D sky130_fd_sc_hd__mux2_1
XFILLER_147_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08083_ _10134_/A0 _10867_/Q _08083_/S vssd1 vssd1 vccd1 vccd1 _08084_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05295_ _11128_/Q _11127_/Q _05393_/S vssd1 vssd1 vccd1 vccd1 _05296_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07034_ _07034_/A _07107_/B vssd1 vssd1 vccd1 vccd1 _07034_/X sky130_fd_sc_hd__and2_1
XFILLER_88_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_124_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11698_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ _11345_/Q _08989_/B vssd1 vssd1 vccd1 vccd1 _08985_/X sky130_fd_sc_hd__or2_1
XFILLER_57_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07936_ _07936_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _10785_/D sky130_fd_sc_hd__or2_1
XFILLER_116_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07867_ _10752_/Q _07883_/B vssd1 vssd1 vccd1 vccd1 _07867_/X sky130_fd_sc_hd__or2_1
X_09606_ _10625_/Q _09947_/A2 _09568_/D _10380_/Q vssd1 vssd1 vccd1 vccd1 _09606_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06818_ _10374_/Q _07203_/A _06858_/B1 _10521_/Q vssd1 vssd1 vccd1 vccd1 _06818_/X
+ sky130_fd_sc_hd__o22a_1
X_07798_ _07916_/A _07798_/B vssd1 vssd1 vccd1 vccd1 _10706_/D sky130_fd_sc_hd__or2_1
X_09537_ _09525_/A _09528_/B _09516_/Y _09536_/X _09825_/A vssd1 vssd1 vccd1 vccd1
+ _11623_/D sky130_fd_sc_hd__o311a_1
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06749_ _10762_/Q _06861_/B _06877_/B1 _10574_/Q vssd1 vssd1 vccd1 vccd1 _06749_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09468_ _09441_/A input24/X _09441_/Y input33/X _09467_/X vssd1 vssd1 vccd1 vccd1
+ _09468_/X sky130_fd_sc_hd__a221o_1
XFILLER_19_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08419_ _09237_/A0 _08414_/S _08418_/X _07003_/B vssd1 vssd1 vccd1 vccd1 _11050_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09399_ _10080_/A0 _11565_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _11565_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11430_ _11431_/CLK _11430_/D vssd1 vssd1 vccd1 vccd1 _11430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11361_ _11811_/CLK _11361_/D vssd1 vssd1 vccd1 vccd1 _11361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10312_ _11308_/CLK _10312_/D vssd1 vssd1 vccd1 vccd1 _10312_/Q sky130_fd_sc_hd__dfxtp_2
X_11292_ _11332_/CLK _11292_/D vssd1 vssd1 vccd1 vccd1 _11292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10243_ _11474_/CLK _10243_/D vssd1 vssd1 vccd1 vccd1 _10243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10174_ _11799_/Q _10176_/B vssd1 vssd1 vccd1 vccd1 _10174_/X sky130_fd_sc_hd__or2_1
XFILLER_105_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11628_ _11628_/CLK _11628_/D vssd1 vssd1 vccd1 vccd1 _11628_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11559_ _11758_/CLK _11559_/D vssd1 vssd1 vccd1 vccd1 _11559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05080_ _11602_/Q vssd1 vssd1 vccd1 vccd1 _09477_/A sky130_fd_sc_hd__clkinv_2
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6__f_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_6__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08770_ _09364_/A1 _11241_/Q _08792_/S vssd1 vssd1 vccd1 vccd1 _08771_/B sky130_fd_sc_hd__mux2_1
X_05982_ _10268_/Q _06858_/B1 _05980_/X _05981_/X vssd1 vssd1 vccd1 vccd1 _05982_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07721_ _09214_/A _07755_/A2 _07720_/X _07868_/C1 vssd1 vssd1 vccd1 vccd1 _10661_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07652_ _08440_/B2 _10616_/Q _07655_/S vssd1 vssd1 vccd1 vccd1 _10616_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06603_ _10778_/Q _06646_/A2 _09131_/A _10667_/Q vssd1 vssd1 vccd1 vccd1 _06603_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07583_ _07034_/A _10575_/Q _07593_/S vssd1 vssd1 vccd1 vccd1 _07584_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09322_ _10080_/A0 _11515_/Q _09324_/S vssd1 vssd1 vccd1 vccd1 _11515_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06534_ _06663_/A _10234_/Q vssd1 vssd1 vccd1 vccd1 _06535_/B sky130_fd_sc_hd__and2_1
XFILLER_0_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09253_ _11479_/Q _09249_/X _09252_/X vssd1 vssd1 vccd1 vccd1 _11479_/D sky130_fd_sc_hd__a21o_1
X_06465_ _10444_/Q _06634_/B1 _06731_/B1 _11078_/Q _11869_/A vssd1 vssd1 vccd1 vccd1
+ _06465_/X sky130_fd_sc_hd__o221a_1
XFILLER_18_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05416_ _10420_/Q _10419_/Q _05416_/S vssd1 vssd1 vccd1 vccd1 _05417_/D sky130_fd_sc_hd__mux2_1
X_08204_ _09393_/A0 _08225_/S _08203_/X _08351_/C1 vssd1 vssd1 vccd1 vccd1 _10936_/D
+ sky130_fd_sc_hd__o211a_1
X_09184_ input101/X _11437_/Q _09184_/S vssd1 vssd1 vccd1 vccd1 _09184_/X sky130_fd_sc_hd__mux2_1
X_06396_ _11082_/Q _08469_/B _06395_/X _06642_/C1 vssd1 vssd1 vccd1 vccd1 _06396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08135_ _08839_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _10893_/D sky130_fd_sc_hd__or2_1
XFILLER_88_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05347_ _11308_/Q _11307_/Q _05382_/S vssd1 vssd1 vccd1 vccd1 _05354_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08066_ _07107_/A _08427_/B _08065_/X _08351_/C1 vssd1 vssd1 vccd1 vccd1 _10858_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05278_ _10821_/Q _10820_/Q _05399_/S vssd1 vssd1 vccd1 vccd1 _05280_/C sky130_fd_sc_hd__mux2_1
XFILLER_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07017_ _10269_/Q _07016_/X _07038_/S vssd1 vssd1 vccd1 vccd1 _10269_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08968_ _11336_/Q _10118_/A0 _08970_/S vssd1 vssd1 vccd1 vccd1 _11336_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07919_ _08935_/A1 _10777_/Q _09221_/C vssd1 vssd1 vccd1 vccd1 _07920_/B sky130_fd_sc_hd__mux2_1
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08899_ _11308_/Q _07309_/X _08901_/S vssd1 vssd1 vccd1 vccd1 _11308_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10930_ _10932_/CLK _10930_/D vssd1 vssd1 vccd1 vccd1 _10930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_92_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11465_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11633_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10861_ _11235_/CLK _10861_/D vssd1 vssd1 vccd1 vccd1 _10861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10792_ _11235_/CLK _10792_/D vssd1 vssd1 vccd1 vccd1 _10792_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11413_ _11792_/CLK _11413_/D vssd1 vssd1 vccd1 vccd1 _11413_/Q sky130_fd_sc_hd__dfxtp_1
X_11344_ _11497_/CLK _11344_/D vssd1 vssd1 vccd1 vccd1 _11344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _11601_/CLK _11275_/D vssd1 vssd1 vccd1 vccd1 _11275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10226_ _10981_/CLK _10226_/D vssd1 vssd1 vccd1 vccd1 _10226_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10157_ _11791_/Q _10137_/X _10156_/X vssd1 vssd1 vccd1 vccd1 _11791_/D sky130_fd_sc_hd__a21o_1
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10088_ _10088_/A1 _10104_/B _10156_/B1 vssd1 vssd1 vccd1 vccd1 _10088_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06250_ _11040_/Q _06735_/A2 _06246_/X _06249_/X vssd1 vssd1 vccd1 vccd1 _06250_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05201_ _05471_/A _08380_/A _05197_/Y _05198_/Y _05200_/Y vssd1 vssd1 vccd1 vccd1
+ _05204_/B sky130_fd_sc_hd__o2111a_1
XFILLER_106_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06181_ _11729_/Q _10061_/A _09347_/A _11534_/Q vssd1 vssd1 vccd1 vccd1 _06181_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_89_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05132_ _10934_/Q _10933_/Q _05399_/S vssd1 vssd1 vccd1 vccd1 _05134_/C sky130_fd_sc_hd__mux2_1
XFILLER_85_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09940_ _11661_/Q _09770_/S _09937_/X _09939_/X vssd1 vssd1 vccd1 vccd1 _11661_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout906 _05093_/Y vssd1 vssd1 vccd1 vccd1 _06450_/A sky130_fd_sc_hd__buf_4
Xfanout917 _06297_/C1 vssd1 vssd1 vccd1 vccd1 _07689_/B sky130_fd_sc_hd__buf_8
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _11399_/Q _09871_/A2 _09565_/D _10573_/Q vssd1 vssd1 vccd1 vccd1 _09871_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout928 _10182_/A0 vssd1 vssd1 vccd1 vccd1 _09393_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 input97/X vssd1 vssd1 vccd1 vccd1 _08893_/A1 sky130_fd_sc_hd__buf_12
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _09396_/A0 _11269_/Q _08838_/S vssd1 vssd1 vccd1 vccd1 _08823_/B sky130_fd_sc_hd__mux2_1
XFILLER_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08753_ _07007_/A _08760_/S _08752_/X _08753_/C1 vssd1 vssd1 vccd1 vccd1 _11233_/D
+ sky130_fd_sc_hd__o211a_1
X_05965_ _11726_/Q _10061_/A _09347_/A _11531_/Q vssd1 vssd1 vccd1 vccd1 _05965_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07704_ _10652_/Q _07693_/Y _07697_/Y _07316_/X vssd1 vssd1 vccd1 vccd1 _10652_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05896_ _05892_/X _05893_/X _05895_/X _07297_/A vssd1 vssd1 vccd1 vccd1 _05896_/X
+ sky130_fd_sc_hd__a31o_2
X_08684_ _08684_/A _08684_/B vssd1 vssd1 vccd1 vccd1 _11196_/D sky130_fd_sc_hd__or2_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07635_ _10604_/Q _07013_/X _07637_/S vssd1 vssd1 vccd1 vccd1 _10604_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07566_ _07918_/A _07566_/B vssd1 vssd1 vccd1 vccd1 _10566_/D sky130_fd_sc_hd__or2_1
XFILLER_146_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09305_ _10171_/A1 _09293_/X _09304_/X _09995_/C1 vssd1 vssd1 vccd1 vccd1 _11503_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06517_ _11435_/Q _06645_/A2 _06648_/A2 _10807_/Q vssd1 vssd1 vccd1 vccd1 _06517_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07497_ _10533_/Q _07537_/B vssd1 vssd1 vccd1 vccd1 _07497_/X sky130_fd_sc_hd__or2_1
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09236_ _11469_/Q _09227_/Y _09228_/Y _07026_/X vssd1 vssd1 vccd1 vccd1 _11469_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_155_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06448_ _11871_/A _06442_/X _06447_/X _06576_/A vssd1 vssd1 vccd1 vccd1 _06448_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09167_ _11428_/Q _09171_/B vssd1 vssd1 vccd1 vccd1 _09167_/X sky130_fd_sc_hd__or2_1
X_06379_ _11198_/Q _06736_/A2 _05789_/Y _06378_/X vssd1 vssd1 vccd1 vccd1 _06379_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08118_ _10886_/Q _08818_/A1 _08120_/S vssd1 vssd1 vccd1 vccd1 _08119_/B sky130_fd_sc_hd__mux2_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ _11396_/Q _09082_/X _09097_/X vssd1 vssd1 vccd1 vccd1 _11396_/D sky130_fd_sc_hd__a21o_1
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08049_ _10851_/Q _08818_/A1 _08051_/S vssd1 vssd1 vccd1 vccd1 _08050_/B sky130_fd_sc_hd__mux2_1
XFILLER_150_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11060_ _11269_/CLK _11060_/D vssd1 vssd1 vccd1 vccd1 _11060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10011_ _07303_/A _11696_/Q _10025_/S vssd1 vssd1 vccd1 vccd1 _10012_/B sky130_fd_sc_hd__mux2_1
XFILLER_103_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ _11220_/CLK _10913_/D vssd1 vssd1 vccd1 vccd1 _10913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10844_ _11224_/CLK _10844_/D vssd1 vssd1 vccd1 vccd1 _10844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10775_ _11472_/CLK _10775_/D vssd1 vssd1 vccd1 vccd1 _10775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11327_ _11329_/CLK _11327_/D vssd1 vssd1 vccd1 vccd1 _11327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11258_ _11572_/CLK _11258_/D vssd1 vssd1 vccd1 vccd1 _11258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10209_ _11808_/CLK _10209_/D vssd1 vssd1 vccd1 vccd1 _10209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11189_ _11325_/CLK _11189_/D vssd1 vssd1 vccd1 vccd1 _11189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05750_ _05751_/A _11868_/A _11867_/A vssd1 vssd1 vccd1 vccd1 _05750_/Y sky130_fd_sc_hd__nor3b_4
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05681_ _11169_/Q _05543_/Y _05597_/Y _11159_/Q vssd1 vssd1 vccd1 vccd1 _05681_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07420_ _07420_/A _07420_/B vssd1 vssd1 vccd1 vccd1 _10486_/D sky130_fd_sc_hd__or2_1
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07351_ _08821_/A _07351_/B vssd1 vssd1 vccd1 vccd1 _10446_/D sky130_fd_sc_hd__and2_1
XFILLER_17_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06302_ _11456_/Q _06862_/A2 _07853_/A _10752_/Q vssd1 vssd1 vccd1 vccd1 _06302_/X
+ sky130_fd_sc_hd__o22a_1
X_07282_ _07922_/A _07282_/B vssd1 vssd1 vccd1 vccd1 _10409_/D sky130_fd_sc_hd__or2_1
XFILLER_137_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06233_ _06224_/X _06226_/X _06227_/X _07690_/A vssd1 vssd1 vccd1 vccd1 _06233_/X
+ sky130_fd_sc_hd__a31o_4
X_09021_ _11361_/Q _09035_/B vssd1 vssd1 vccd1 vccd1 _09021_/X sky130_fd_sc_hd__or2_1
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06164_ _10639_/Q _06538_/B1 _06504_/B1 _10952_/Q vssd1 vssd1 vccd1 vccd1 _06164_/X
+ sky130_fd_sc_hd__o22a_1
X_05115_ _11178_/Q _10303_/Q _05392_/S vssd1 vssd1 vccd1 vccd1 _05118_/B sky130_fd_sc_hd__mux2_1
XFILLER_89_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06095_ _11728_/Q _08200_/A _09347_/A _11533_/Q vssd1 vssd1 vccd1 vccd1 _06095_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_104_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09923_ _10490_/Q _09570_/A _09565_/A _10487_/Q vssd1 vssd1 vccd1 vccd1 _09923_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout703 _05380_/S vssd1 vssd1 vccd1 vccd1 _05418_/S sky130_fd_sc_hd__buf_6
Xfanout714 _06556_/B1 vssd1 vssd1 vccd1 vccd1 _08647_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout725 fanout726/X vssd1 vssd1 vccd1 vccd1 _06540_/B1 sky130_fd_sc_hd__buf_4
Xfanout736 _08765_/A vssd1 vssd1 vccd1 vccd1 _06716_/B1 sky130_fd_sc_hd__clkbuf_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ _10701_/Q _09873_/A2 _09873_/B1 _10707_/Q _09853_/X vssd1 vssd1 vccd1 vccd1
+ _09861_/A sky130_fd_sc_hd__a221o_1
Xfanout747 _08472_/A vssd1 vssd1 vccd1 vccd1 _06629_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout758 _06674_/A2 vssd1 vssd1 vccd1 vccd1 _06875_/B1 sky130_fd_sc_hd__buf_6
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout769 _10119_/A vssd1 vssd1 vccd1 vccd1 _05865_/B sky130_fd_sc_hd__buf_6
XFILLER_85_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _08947_/A1 _08802_/S _08804_/X _08947_/C1 vssd1 vssd1 vccd1 vccd1 _11258_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09785_ _11648_/Q _09404_/Y _09784_/X _09681_/B vssd1 vssd1 vccd1 vccd1 _09785_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06997_ _06997_/A _07151_/B _07151_/C _07151_/D vssd1 vssd1 vccd1 vccd1 _06997_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08736_ _07021_/A _11225_/Q _08748_/S vssd1 vssd1 vccd1 vccd1 _08737_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05948_ _06535_/A _05886_/X _05947_/X _06664_/C1 vssd1 vssd1 vccd1 vccd1 _05950_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 fanout755/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_118 _09081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _10177_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ _08668_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08705_/B sky130_fd_sc_hd__nor2_4
XFILLER_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05879_ _11088_/Q _06629_/B1 _05877_/X _05878_/X vssd1 vssd1 vccd1 vccd1 _05879_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07618_ _10593_/Q _07613_/Y _07614_/Y _07617_/X vssd1 vssd1 vccd1 vccd1 _10593_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08598_ _09114_/A1 _08623_/S _08597_/X _08947_/C1 vssd1 vssd1 vccd1 vccd1 _11153_/D
+ sky130_fd_sc_hd__o211a_1
X_07549_ _10017_/A0 _10558_/Q _07589_/S vssd1 vssd1 vccd1 vccd1 _07550_/B sky130_fd_sc_hd__mux2_1
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10560_ _10773_/CLK _10560_/D vssd1 vssd1 vccd1 vccd1 _10560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ _07441_/A _09218_/X _09241_/B1 vssd1 vssd1 vccd1 vccd1 _11458_/D sky130_fd_sc_hd__o21a_1
XFILLER_108_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ _11706_/CLK _10491_/D vssd1 vssd1 vccd1 vccd1 _10491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11112_ _11319_/CLK _11112_/D vssd1 vssd1 vccd1 vccd1 _11112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11043_ _11575_/CLK _11043_/D vssd1 vssd1 vccd1 vccd1 _11043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10827_ _10939_/CLK _10827_/D vssd1 vssd1 vccd1 vccd1 _10827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10758_ _11470_/CLK _10758_/D vssd1 vssd1 vccd1 vccd1 _10758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10689_ _10735_/CLK _10689_/D vssd1 vssd1 vccd1 vccd1 _10689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06920_ _10105_/A1 _06922_/B _08664_/A vssd1 vssd1 vccd1 vccd1 _06920_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06851_ _06841_/X _06842_/X _06845_/X _06850_/X vssd1 vssd1 vccd1 vccd1 _06851_/X
+ sky130_fd_sc_hd__a31o_1
X_05802_ _11181_/Q _07190_/A _05800_/X _05801_/X vssd1 vssd1 vccd1 vccd1 _05802_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_1363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09570_ _09570_/A _09570_/B vssd1 vssd1 vccd1 vccd1 _09574_/A sky130_fd_sc_hd__or2_1
X_06782_ _06853_/A1 _10244_/Q _06852_/A3 _06743_/X _06781_/X vssd1 vssd1 vccd1 vccd1
+ _06782_/X sky130_fd_sc_hd__a32o_1
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08521_ _11110_/Q _08545_/B vssd1 vssd1 vccd1 vccd1 _08521_/X sky130_fd_sc_hd__or2_1
X_05733_ _05819_/A _06892_/B vssd1 vssd1 vccd1 vccd1 _06743_/A sky130_fd_sc_hd__nor2_8
XFILLER_70_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08452_ _11073_/Q _08459_/S _07628_/S _07229_/B vssd1 vssd1 vccd1 vccd1 _11073_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_50_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05664_ _11255_/Q _05579_/Y _05597_/Y _11246_/Q vssd1 vssd1 vccd1 vccd1 _05664_/X
+ sky130_fd_sc_hd__a22o_1
X_07403_ _10017_/A0 _10478_/Q _07425_/S vssd1 vssd1 vccd1 vccd1 _07404_/B sky130_fd_sc_hd__mux2_1
X_05595_ _05619_/A1 _11487_/Q _11483_/Q _05619_/B2 _05593_/X vssd1 vssd1 vccd1 vccd1
+ _05595_/X sky130_fd_sc_hd__a221o_1
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08383_ _08383_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08383_/X sky130_fd_sc_hd__or2_4
XFILLER_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07334_ _10433_/Q _07322_/Y _07326_/Y _07333_/X vssd1 vssd1 vccd1 vccd1 _10433_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07265_ _09214_/A _10401_/Q _09187_/S vssd1 vssd1 vccd1 vccd1 _07266_/B sky130_fd_sc_hd__mux2_1
X_09004_ _10185_/A0 _08994_/X _09003_/X _09036_/C1 vssd1 vssd1 vccd1 vccd1 _11353_/D
+ sky130_fd_sc_hd__o211a_1
X_06216_ _11545_/Q _06219_/A2 _06214_/X _06215_/X vssd1 vssd1 vccd1 vccd1 _06216_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07196_ _07141_/B _07195_/X _07318_/A vssd1 vssd1 vccd1 vccd1 _10358_/D sky130_fd_sc_hd__a21o_1
XFILLER_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06147_ _11183_/Q _08650_/A _06639_/B1 _10814_/Q vssd1 vssd1 vccd1 vccd1 _06151_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06078_ _07082_/A _06076_/X _06077_/X _06075_/X _05816_/A vssd1 vssd1 vccd1 vccd1
+ _06078_/X sky130_fd_sc_hd__a221o_1
XFILLER_105_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout500 _09048_/C1 vssd1 vssd1 vccd1 vccd1 _08943_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout511 _08819_/A vssd1 vssd1 vccd1 vccd1 _08810_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09906_ _11706_/Q _09947_/A2 _09572_/B _11718_/Q _09905_/X vssd1 vssd1 vccd1 vccd1
+ _09907_/D sky130_fd_sc_hd__a221o_1
Xfanout522 _07659_/A vssd1 vssd1 vccd1 vccd1 _07664_/A sky130_fd_sc_hd__buf_4
Xfanout533 fanout536/X vssd1 vssd1 vccd1 vccd1 _10150_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout544 _07918_/A vssd1 vssd1 vccd1 vccd1 _07934_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout555 _06898_/Y vssd1 vssd1 vccd1 vccd1 fanout555/X sky130_fd_sc_hd__buf_6
XFILLER_63_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout566 _06898_/Y vssd1 vssd1 vccd1 vccd1 _08773_/A sky130_fd_sc_hd__buf_4
Xfanout577 fanout578/X vssd1 vssd1 vccd1 vccd1 _09129_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_112_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _10775_/Q _09573_/A _09953_/B1 _11463_/Q _09836_/X vssd1 vssd1 vccd1 vccd1
+ _09842_/B sky130_fd_sc_hd__a221o_1
XFILLER_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout588 _05734_/X vssd1 vssd1 vccd1 vccd1 _06852_/A3 sky130_fd_sc_hd__buf_6
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout599 _05789_/Y vssd1 vssd1 vccd1 vccd1 _06718_/C1 sky130_fd_sc_hd__buf_6
XFILLER_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09768_ _09497_/A _09722_/Y _09758_/Y _06969_/X vssd1 vssd1 vccd1 vccd1 _09768_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _08810_/A _08719_/B vssd1 vssd1 vccd1 vccd1 _11215_/D sky130_fd_sc_hd__or2_1
XFILLER_26_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09699_ _09703_/A _09699_/B vssd1 vssd1 vccd1 vccd1 _11640_/D sky130_fd_sc_hd__or2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11735_/CLK _11730_/D vssd1 vssd1 vccd1 vccd1 _11730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11661_/CLK _11661_/D vssd1 vssd1 vccd1 vccd1 _11661_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10612_ _11777_/CLK _10612_/D vssd1 vssd1 vccd1 vccd1 _10612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11592_ _11604_/CLK _11592_/D vssd1 vssd1 vccd1 vccd1 _11592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10543_ _10782_/CLK _10543_/D vssd1 vssd1 vccd1 vccd1 _10543_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_109_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10474_ _11706_/CLK _10474_/D vssd1 vssd1 vccd1 vccd1 _10474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11026_ _11270_/CLK _11026_/D vssd1 vssd1 vccd1 vccd1 _11026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05380_ _10617_/Q _10616_/Q _05380_/S vssd1 vssd1 vccd1 vccd1 _05384_/A sky130_fd_sc_hd__mux2_1
XANTENNA_18 _06387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 _07008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07050_ _10281_/Q _07047_/B _07491_/S _07005_/A vssd1 vssd1 vccd1 vccd1 _10281_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06001_ _10823_/Q _06415_/A2 _06453_/B1 _10988_/Q vssd1 vssd1 vccd1 vccd1 _06001_/X
+ sky130_fd_sc_hd__o22a_1
Xoutput125 _05704_/X vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_4
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput136 _11616_/Q vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_4
Xoutput147 _11570_/Q vssd1 vssd1 vccd1 vccd1 ram_addr[1] sky130_fd_sc_hd__buf_4
Xoutput158 _11578_/Q vssd1 vssd1 vccd1 vccd1 rom_addr[0] sky130_fd_sc_hd__buf_4
XFILLER_115_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput169 _11867_/X vssd1 vssd1 vccd1 vccd1 wb_rom_adrb[1] sky130_fd_sc_hd__buf_4
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07952_ _10794_/Q _07942_/Y _07943_/Y _07335_/X vssd1 vssd1 vccd1 vccd1 _10794_/D
+ sky130_fd_sc_hd__o22a_1
X_06903_ _06903_/A _10180_/C _10137_/B vssd1 vssd1 vccd1 vccd1 _06903_/X sky130_fd_sc_hd__or3_4
X_07883_ _10760_/Q _07883_/B vssd1 vssd1 vccd1 vccd1 _07883_/X sky130_fd_sc_hd__or2_1
X_09622_ _10719_/Q _09568_/B _09571_/C _10733_/Q vssd1 vssd1 vccd1 vccd1 _09622_/X
+ sky130_fd_sc_hd__a22o_1
X_06834_ _10766_/Q _07854_/A _06875_/B1 _10679_/Q vssd1 vssd1 vccd1 vccd1 _06834_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09553_ _09553_/A _09668_/B _09668_/C vssd1 vssd1 vccd1 vccd1 _09673_/B sky130_fd_sc_hd__nor3_4
X_06765_ _10713_/Q _07777_/A _06877_/B1 _10575_/Q _06764_/X vssd1 vssd1 vccd1 vccd1
+ _06765_/X sky130_fd_sc_hd__o221a_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08504_ _08665_/A _08501_/S _08503_/X _08662_/C1 vssd1 vssd1 vccd1 vccd1 _11102_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05716_ _05716_/A _05716_/B _05716_/C _05716_/D vssd1 vssd1 vccd1 vccd1 _05716_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_110_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09484_ _09515_/B _09515_/C vssd1 vssd1 vccd1 vccd1 _09504_/B sky130_fd_sc_hd__nor2_1
X_06696_ _11050_/Q _06696_/A2 _08245_/A _10972_/Q vssd1 vssd1 vccd1 vccd1 _06696_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08435_ _11060_/Q _08424_/Y _08427_/Y _07019_/X vssd1 vssd1 vccd1 vccd1 _11060_/D
+ sky130_fd_sc_hd__a22o_1
X_05647_ _11303_/Q _05591_/Y _05633_/Y _11286_/Q vssd1 vssd1 vccd1 vccd1 _05655_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08366_ _11025_/Q _08438_/B vssd1 vssd1 vccd1 vccd1 _08366_/X sky130_fd_sc_hd__or2_1
X_05578_ _05626_/A2 _11365_/Q _11360_/Q _05630_/B1 _05577_/X vssd1 vssd1 vccd1 vccd1
+ _05579_/B sky130_fd_sc_hd__a221o_4
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07317_ _10425_/Q _07301_/Y _07306_/Y _07316_/X vssd1 vssd1 vccd1 vccd1 _10425_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08297_ _10983_/Q _07100_/X _08298_/S vssd1 vssd1 vccd1 vccd1 _10983_/D sky130_fd_sc_hd__mux2_1
X_07248_ _10051_/A1 _07141_/B _07318_/A vssd1 vssd1 vccd1 vccd1 _07248_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_46_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11791_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_106_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07179_ _10047_/A1 _09240_/S _07178_/X _07932_/C1 vssd1 vssd1 vccd1 vccd1 _10350_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10190_ _10190_/A0 _11811_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _11811_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout330 _07172_/S vssd1 vssd1 vccd1 vccd1 _09243_/C sky130_fd_sc_hd__buf_6
Xfanout341 _08907_/B vssd1 vssd1 vccd1 vccd1 _08906_/B sky130_fd_sc_hd__buf_12
Xfanout352 _07643_/C vssd1 vssd1 vccd1 vccd1 _08471_/B sky130_fd_sc_hd__buf_6
Xfanout363 _07335_/B vssd1 vssd1 vccd1 vccd1 _08817_/B2 sky130_fd_sc_hd__buf_8
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout374 _08322_/A vssd1 vssd1 vccd1 vccd1 _07318_/A sky130_fd_sc_hd__buf_6
Xfanout385 _07614_/A vssd1 vssd1 vccd1 vccd1 _09229_/A sky130_fd_sc_hd__buf_12
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout396 _07003_/Y vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__buf_12
XFILLER_115_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11713_/CLK _11713_/D vssd1 vssd1 vccd1 vccd1 _11713_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11644_/CLK _11644_/D vssd1 vssd1 vccd1 vccd1 _11644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11575_ _11575_/CLK _11575_/D vssd1 vssd1 vccd1 vccd1 _11575_/Q sky130_fd_sc_hd__dfxtp_4
Xinput16 rom_value[15] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_2
Xinput27 rom_value[25] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput38 rom_value[6] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10526_ _11706_/CLK _10526_/D vssd1 vssd1 vccd1 vccd1 _10526_/Q sky130_fd_sc_hd__dfxtp_2
Xinput49 wb_rom_val[16] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_4
XFILLER_156_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10457_ _11308_/CLK _10457_/D vssd1 vssd1 vccd1 vccd1 _10457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10388_ _11711_/CLK _10388_/D vssd1 vssd1 vccd1 vccd1 _10388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_5__f_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_5__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11009_ _11067_/CLK _11009_/D vssd1 vssd1 vccd1 vccd1 _11009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06550_ _10740_/Q _06634_/B1 _06731_/B1 _10599_/Q _06550_/C1 vssd1 vssd1 vccd1 vccd1
+ _06550_/X sky130_fd_sc_hd__o221a_1
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05501_ _10246_/Q input58/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05501_/X sky130_fd_sc_hd__mux2_2
X_06481_ _10367_/Q _09358_/A _09976_/A _10512_/Q _07151_/A vssd1 vssd1 vccd1 vccd1
+ _06481_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08220_ _08492_/A _08220_/B vssd1 vssd1 vccd1 vccd1 _10944_/D sky130_fd_sc_hd__or2_1
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05432_ _10651_/Q _10650_/Q _05432_/S vssd1 vssd1 vccd1 vccd1 _05433_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05363_ _10986_/Q _10985_/Q _05427_/S vssd1 vssd1 vccd1 vccd1 _05367_/A sky130_fd_sc_hd__mux2_2
X_08151_ _10182_/A0 _08162_/S _08150_/X _08753_/C1 vssd1 vssd1 vccd1 vccd1 _10901_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07102_ _07617_/A _07318_/B vssd1 vssd1 vccd1 vccd1 _07102_/X sky130_fd_sc_hd__or2_2
X_05294_ _11126_/Q _11125_/Q _05396_/S vssd1 vssd1 vccd1 vccd1 _05296_/C sky130_fd_sc_hd__mux2_1
X_08082_ _07061_/A _08083_/S _08081_/X _08753_/C1 vssd1 vssd1 vccd1 vccd1 _10866_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07033_ _09229_/A _07033_/B vssd1 vssd1 vccd1 vccd1 _10275_/D sky130_fd_sc_hd__and2_1
XFILLER_106_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08984_ _11344_/Q _08972_/X _08983_/X vssd1 vssd1 vccd1 vccd1 _11344_/D sky130_fd_sc_hd__a21o_1
XFILLER_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07935_ input103/X _10785_/Q _09206_/B vssd1 vssd1 vccd1 vccd1 _07936_/B sky130_fd_sc_hd__mux2_1
XFILLER_60_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07866_ _10023_/A0 _07871_/S _07865_/X _07866_/C1 vssd1 vssd1 vccd1 vccd1 _10751_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09605_ _10390_/Q _09567_/B _09570_/B _10389_/Q vssd1 vssd1 vccd1 vccd1 _09605_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06817_ _11473_/Q _07153_/A _06816_/X _06878_/C1 vssd1 vssd1 vccd1 vccd1 _06817_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07797_ _08931_/A1 _10706_/Q _09193_/B vssd1 vssd1 vccd1 vccd1 _07798_/B sky130_fd_sc_hd__mux2_1
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09536_ _09492_/B _09489_/C _09516_/A _11623_/Q vssd1 vssd1 vccd1 vccd1 _09536_/X
+ sky130_fd_sc_hd__a31o_1
X_06748_ _10712_/Q _06748_/A2 _07440_/A _10547_/Q vssd1 vssd1 vccd1 vccd1 _06748_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_145_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09467_ _09441_/A input15/X _09441_/B vssd1 vssd1 vccd1 vccd1 _09467_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06679_ _11329_/Q _06738_/A2 _06739_/A2 _11301_/Q _05789_/Y vssd1 vssd1 vccd1 vccd1
+ _06679_/X sky130_fd_sc_hd__o221a_1
XFILLER_145_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08418_ _11050_/Q _08422_/B vssd1 vssd1 vccd1 vccd1 _08418_/X sky130_fd_sc_hd__or2_1
X_09398_ _10115_/A0 _11564_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _11564_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08349_ _08835_/A _08349_/B vssd1 vssd1 vccd1 vccd1 _11017_/D sky130_fd_sc_hd__or2_1
XFILLER_123_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _11607_/CLK _11360_/D vssd1 vssd1 vccd1 vccd1 _11360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10311_ _10798_/CLK _10311_/D vssd1 vssd1 vccd1 vccd1 _10311_/Q sky130_fd_sc_hd__dfxtp_1
X_11291_ _11291_/CLK _11291_/D vssd1 vssd1 vccd1 vccd1 _11291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10242_ _11712_/CLK _10242_/D vssd1 vssd1 vccd1 vccd1 _10242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10173_ _11798_/Q _10159_/X _10172_/X vssd1 vssd1 vccd1 vccd1 _11798_/D sky130_fd_sc_hd__a21o_1
XFILLER_105_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11627_ _11657_/CLK _11627_/D vssd1 vssd1 vccd1 vccd1 _11627_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11558_ _11675_/CLK _11558_/D vssd1 vssd1 vccd1 vccd1 _11558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10509_ _11702_/CLK _10509_/D vssd1 vssd1 vccd1 vccd1 _10509_/Q sky130_fd_sc_hd__dfxtp_1
X_11489_ _11497_/CLK _11489_/D vssd1 vssd1 vccd1 vccd1 _11489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05981_ _10477_/Q _06872_/A2 _10009_/A _11743_/Q _06849_/C1 vssd1 vssd1 vccd1 vccd1
+ _05981_/X sky130_fd_sc_hd__o221a_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07720_ _10661_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07720_/X sky130_fd_sc_hd__or2_1
X_07651_ _10615_/Q _08901_/A1 _07651_/S vssd1 vssd1 vccd1 vccd1 _10615_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06602_ _11436_/Q _06645_/A2 _08971_/A _10568_/Q vssd1 vssd1 vccd1 vccd1 _06602_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07582_ _07930_/A _07582_/B vssd1 vssd1 vccd1 vccd1 _10574_/D sky130_fd_sc_hd__or2_1
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09321_ _10115_/A0 _11514_/Q _09324_/S vssd1 vssd1 vccd1 vccd1 _11514_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06533_ _11871_/A _06527_/X _06532_/X _07081_/A _06516_/X vssd1 vssd1 vccd1 vccd1
+ _06533_/X sky130_fd_sc_hd__a32o_1
XFILLER_80_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _10182_/A0 _09266_/B _08761_/A vssd1 vssd1 vccd1 vccd1 _09252_/X sky130_fd_sc_hd__a21o_1
XFILLER_90_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06464_ _10920_/Q _06591_/A2 _06126_/B _10745_/Q vssd1 vssd1 vccd1 vccd1 _06467_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_142_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08203_ _10936_/Q _08902_/C vssd1 vssd1 vccd1 vccd1 _08203_/X sky130_fd_sc_hd__or2_1
X_05415_ _11234_/Q _11233_/Q _06939_/A vssd1 vssd1 vccd1 vccd1 _05417_/C sky130_fd_sc_hd__mux2_1
X_09183_ _07441_/A _09182_/X _09241_/B1 vssd1 vssd1 vccd1 vccd1 _11436_/D sky130_fd_sc_hd__o21a_1
X_06395_ _10847_/Q _06643_/A2 _08650_/A _11226_/Q _06394_/X vssd1 vssd1 vccd1 vccd1
+ _06395_/X sky130_fd_sc_hd__o221a_1
XFILLER_147_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08134_ _09323_/A0 _10893_/Q _08146_/S vssd1 vssd1 vccd1 vccd1 _08135_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05346_ _05346_/A _05346_/B vssd1 vssd1 vccd1 vccd1 _05346_/Y sky130_fd_sc_hd__nor2_8
XFILLER_105_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08065_ _10858_/Q _08426_/B vssd1 vssd1 vccd1 vccd1 _08065_/X sky130_fd_sc_hd__or2_1
X_05277_ _10819_/Q _10818_/Q _05397_/S vssd1 vssd1 vccd1 vccd1 _05280_/B sky130_fd_sc_hd__mux2_1
X_07016_ _08438_/A _07095_/B vssd1 vssd1 vccd1 vccd1 _07016_/X sky130_fd_sc_hd__or2_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08967_ _11335_/Q _09323_/A0 _08970_/S vssd1 vssd1 vccd1 vccd1 _11335_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07918_ _07918_/A _07918_/B vssd1 vssd1 vccd1 vccd1 _10776_/D sky130_fd_sc_hd__or2_1
XFILLER_56_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08898_ _11307_/Q _07229_/X _08901_/S vssd1 vssd1 vccd1 vccd1 _11307_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07849_ _08440_/B2 _10742_/Q _07852_/S vssd1 vssd1 vccd1 vccd1 _10742_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10860_ _10939_/CLK _10860_/D vssd1 vssd1 vccd1 vccd1 _10860_/Q sky130_fd_sc_hd__dfxtp_1
X_09519_ _09497_/A _09485_/X _09489_/C _11616_/Q vssd1 vssd1 vccd1 vccd1 _09519_/X
+ sky130_fd_sc_hd__a31o_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10791_ _11005_/CLK _10791_/D vssd1 vssd1 vccd1 vccd1 _10791_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_wb_clk_i clkbuf_leaf_69_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11683_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11412_ _11801_/CLK _11412_/D vssd1 vssd1 vccd1 vccd1 _11412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11343_ _11495_/CLK _11343_/D vssd1 vssd1 vccd1 vccd1 _11343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11274_ _11634_/CLK _11274_/D vssd1 vssd1 vccd1 vccd1 _11274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10225_ _11233_/CLK _10225_/D vssd1 vssd1 vccd1 vccd1 _10225_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_106_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10156_ _07057_/A _10154_/B _10156_/B1 vssd1 vssd1 vccd1 vccd1 _10156_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10087_ _10087_/A _10137_/B _10087_/C vssd1 vssd1 vccd1 vccd1 _10087_/X sky130_fd_sc_hd__or3_4
XFILLER_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10989_ _11633_/CLK _10989_/D vssd1 vssd1 vccd1 vccd1 _10989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05200_ _05471_/A _11031_/Q vssd1 vssd1 vccd1 vccd1 _05200_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06180_ _11692_/Q _09998_/A _06924_/A _11739_/Q _06344_/C1 vssd1 vssd1 vccd1 vccd1
+ _06180_/X sky130_fd_sc_hd__o221a_1
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05131_ _10932_/Q _10931_/Q _05397_/S vssd1 vssd1 vccd1 vccd1 _05134_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout907 _05093_/Y vssd1 vssd1 vccd1 vccd1 _06663_/A sky130_fd_sc_hd__clkbuf_4
X_09870_ _11662_/Q _09938_/B vssd1 vssd1 vccd1 vccd1 _09870_/Y sky130_fd_sc_hd__nor2_1
Xfanout918 _06808_/C1 vssd1 vssd1 vccd1 vccd1 _06878_/C1 sky130_fd_sc_hd__buf_6
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 _07002_/A vssd1 vssd1 vccd1 vccd1 _10182_/A0 sky130_fd_sc_hd__buf_6
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08821_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _11268_/D sky130_fd_sc_hd__and2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _11233_/Q _08762_/B vssd1 vssd1 vccd1 vccd1 _08752_/X sky130_fd_sc_hd__or2_1
X_05964_ _11689_/Q _09998_/A _06924_/A _11736_/Q _06344_/C1 vssd1 vssd1 vccd1 vccd1
+ _05964_/X sky130_fd_sc_hd__o221a_1
XFILLER_38_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07703_ _10651_/Q _07694_/Y _07696_/Y _07314_/X vssd1 vssd1 vccd1 vccd1 _10651_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_113_1364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08683_ _08987_/A1 _11196_/Q _08683_/S vssd1 vssd1 vccd1 vccd1 _08684_/B sky130_fd_sc_hd__mux2_1
X_05895_ _11381_/Q _09060_/A _08972_/A _11341_/Q _05894_/X vssd1 vssd1 vccd1 vccd1
+ _05895_/X sky130_fd_sc_hd__o221a_1
XFILLER_66_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07634_ _10603_/Q _07008_/X _07637_/S vssd1 vssd1 vccd1 vccd1 _10603_/D sky130_fd_sc_hd__mux2_1
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07565_ _08846_/A0 _10566_/Q _07593_/S vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__mux2_1
XFILLER_94_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09304_ _11503_/Q _09310_/B vssd1 vssd1 vccd1 vccd1 _09304_/X sky130_fd_sc_hd__or2_1
X_06516_ _06500_/X _06505_/X _06510_/X _06515_/X vssd1 vssd1 vccd1 vccd1 _06516_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07496_ _07043_/X _10532_/Q _07496_/S vssd1 vssd1 vccd1 vccd1 _10532_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09235_ _10043_/A _09234_/X _09243_/B vssd1 vssd1 vccd1 vccd1 _11468_/D sky130_fd_sc_hd__o21a_1
XFILLER_10_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06447_ _11162_/Q _06649_/A2 _06443_/X _06446_/X vssd1 vssd1 vccd1 vccd1 _06447_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_107_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09166_ _10171_/A1 _09154_/X _09165_/X _10175_/C1 vssd1 vssd1 vccd1 vccd1 _11427_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06378_ _11042_/Q _06735_/A2 _08765_/A _11248_/Q _06377_/X vssd1 vssd1 vccd1 vccd1
+ _06378_/X sky130_fd_sc_hd__o221a_1
XFILLER_147_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08117_ _10885_/Q _08120_/S _07642_/S _08817_/B2 vssd1 vssd1 vccd1 vccd1 _10885_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05329_ _05329_/A _05329_/B _05329_/C _05329_/D vssd1 vssd1 vccd1 vccd1 _05335_/A
+ sky130_fd_sc_hd__or4_4
X_09097_ _10023_/A0 _09099_/B _08873_/A vssd1 vssd1 vccd1 vccd1 _09097_/X sky130_fd_sc_hd__a21o_1
X_08048_ _10850_/Q _08051_/S _07365_/Y _08817_/B2 vssd1 vssd1 vccd1 vccd1 _10850_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_150_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10010_ _10010_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _10025_/S sky130_fd_sc_hd__or2_4
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09999_ _09999_/A0 _11686_/Q _10008_/S vssd1 vssd1 vccd1 vccd1 _11686_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10912_ _11779_/CLK _10912_/D vssd1 vssd1 vccd1 vccd1 _10912_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10843_ _11527_/CLK _10843_/D vssd1 vssd1 vccd1 vccd1 _10843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10774_ _11465_/CLK _10774_/D vssd1 vssd1 vccd1 vccd1 _10774_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_13_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11326_ _11330_/CLK _11326_/D vssd1 vssd1 vccd1 vccd1 _11326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11257_ _11291_/CLK _11257_/D vssd1 vssd1 vccd1 vccd1 _11257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10208_ _11810_/CLK _10208_/D vssd1 vssd1 vccd1 vccd1 _10208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11188_ _11607_/CLK _11188_/D vssd1 vssd1 vccd1 vccd1 _11188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10139_ _10181_/A0 _10137_/X _10138_/X _10153_/C1 vssd1 vssd1 vccd1 vccd1 _11782_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05680_ _05680_/A _05680_/B _05680_/C _05680_/D vssd1 vssd1 vccd1 vccd1 _05680_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07350_ _10446_/Q _08647_/A _07350_/S vssd1 vssd1 vccd1 vccd1 _07351_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06301_ _10401_/Q _06804_/B _07540_/A _10562_/Q vssd1 vssd1 vccd1 vccd1 _06301_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_143_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07281_ _07031_/A _10409_/Q _09184_/S vssd1 vssd1 vccd1 vccd1 _07282_/B sky130_fd_sc_hd__mux2_1
XFILLER_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09020_ _11360_/Q _09016_/X _09019_/X vssd1 vssd1 vccd1 vccd1 _11360_/D sky130_fd_sc_hd__a21o_1
X_06232_ _10210_/Q _06351_/A2 _06228_/X _06231_/X vssd1 vssd1 vccd1 vccd1 _06232_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_15_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06163_ _10585_/Q _06454_/A2 _06455_/B1 _10904_/Q vssd1 vssd1 vccd1 vccd1 _06163_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_145_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05114_ _10307_/Q _10306_/Q _05385_/S vssd1 vssd1 vccd1 vccd1 _05118_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06094_ _11671_/Q _09965_/A _08311_/A _10996_/Q vssd1 vssd1 vccd1 vccd1 _06094_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_116_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09922_ _10360_/Q _09571_/C _09572_/D _10482_/Q _09921_/X vssd1 vssd1 vccd1 vccd1
+ _09925_/C sky130_fd_sc_hd__a221o_1
XFILLER_132_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout704 _11594_/Q vssd1 vssd1 vccd1 vccd1 _05380_/S sky130_fd_sc_hd__buf_4
XFILLER_113_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout715 _06556_/B1 vssd1 vssd1 vccd1 vccd1 _08469_/B sky130_fd_sc_hd__buf_6
XFILLER_63_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout726 fanout738/X vssd1 vssd1 vccd1 vccd1 fanout726/X sky130_fd_sc_hd__buf_8
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09853_ _10715_/Q _09872_/A2 _09872_/B1 _10702_/Q vssd1 vssd1 vccd1 vccd1 _09853_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout737 fanout738/X vssd1 vssd1 vccd1 vccd1 _08765_/A sky130_fd_sc_hd__clkbuf_16
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout748 _08472_/A vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__buf_6
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout759 _06674_/A2 vssd1 vssd1 vccd1 vccd1 _07455_/A sky130_fd_sc_hd__buf_6
XFILLER_86_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08804_ _11258_/Q _08804_/B vssd1 vssd1 vccd1 vccd1 _08804_/X sky130_fd_sc_hd__or2_1
X_09784_ _11649_/Q _09771_/Y _09783_/X _09554_/B _09406_/B vssd1 vssd1 vccd1 vccd1
+ _09784_/X sky130_fd_sc_hd__o221a_1
X_06996_ _10106_/A1 _06976_/X _06995_/X _06996_/C1 vssd1 vssd1 vccd1 vccd1 _10265_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08735_ _07052_/A _08742_/S _08734_/X _07107_/B vssd1 vssd1 vccd1 vccd1 _11224_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05947_ _07082_/A _05945_/X _05946_/X _05816_/A vssd1 vssd1 vccd1 vccd1 _05947_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_108 fanout755/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_119 _09216_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _11188_/Q _08663_/S _08665_/X _09036_/C1 vssd1 vssd1 vccd1 vccd1 _11188_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05878_ _10936_/Q _06630_/A2 _06630_/B1 _11012_/Q vssd1 vssd1 vccd1 vccd1 _05878_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_54_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _07617_/A _07617_/B vssd1 vssd1 vccd1 vccd1 _07617_/X sky130_fd_sc_hd__or2_4
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ _11153_/Q _08633_/B vssd1 vssd1 vccd1 vccd1 _08597_/X sky130_fd_sc_hd__or2_1
XFILLER_81_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07548_ _07928_/A _07548_/B vssd1 vssd1 vccd1 vccd1 _10557_/D sky130_fd_sc_hd__or2_1
XFILLER_70_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07479_ _10051_/A1 _10518_/Q _07483_/S vssd1 vssd1 vccd1 vccd1 _07480_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09218_ input101/X _11458_/Q _09218_/S vssd1 vssd1 vccd1 vccd1 _09218_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10490_ _11712_/CLK _10490_/D vssd1 vssd1 vccd1 vccd1 _10490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09149_ _11420_/Q _09149_/B vssd1 vssd1 vccd1 vccd1 _09149_/X sky130_fd_sc_hd__or2_1
XFILLER_33_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11111_ _11428_/CLK _11111_/D vssd1 vssd1 vccd1 vccd1 _11111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11042_ _11319_/CLK _11042_/D vssd1 vssd1 vccd1 vccd1 _11042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10826_ _11601_/CLK _10826_/D vssd1 vssd1 vccd1 vccd1 _10826_/Q sky130_fd_sc_hd__dfxtp_1
X_10757_ _11472_/CLK _10757_/D vssd1 vssd1 vccd1 vccd1 _10757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ _10981_/CLK _10688_/D vssd1 vssd1 vccd1 vccd1 _10688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11309_ _11776_/CLK _11309_/D vssd1 vssd1 vccd1 vccd1 _11309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06850_ _10361_/Q _06872_/A2 _06846_/X _06849_/X vssd1 vssd1 vccd1 vccd1 _06850_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05801_ _10616_/Q _06371_/A2 _07827_/A2 _10975_/Q vssd1 vssd1 vccd1 vccd1 _05801_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_23_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06781_ _06776_/X _06777_/X _06780_/X _06775_/X vssd1 vssd1 vccd1 vccd1 _06781_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_36_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08520_ _08875_/A _08520_/B vssd1 vssd1 vccd1 vccd1 _11109_/D sky130_fd_sc_hd__or2_1
X_05732_ input77/X _10255_/D vssd1 vssd1 vccd1 vccd1 _06892_/B sky130_fd_sc_hd__nand2_8
X_08451_ _11072_/Q _08459_/S _07628_/S _07227_/B vssd1 vssd1 vccd1 vccd1 _11072_/D
+ sky130_fd_sc_hd__o22a_1
X_05663_ _11257_/Q _05591_/Y _05633_/Y _11240_/Q _05662_/X vssd1 vssd1 vccd1 vccd1
+ _05668_/B sky130_fd_sc_hd__a221o_2
XFILLER_23_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07402_ _10050_/A _07402_/B vssd1 vssd1 vccd1 vccd1 _10477_/D sky130_fd_sc_hd__or2_1
X_08382_ _09060_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08422_/B sky130_fd_sc_hd__nor2_8
X_05594_ _05630_/A2 _11481_/Q _11478_/Q _05079_/A _05592_/X vssd1 vssd1 vccd1 vccd1
+ _05597_/A sky130_fd_sc_hd__a221o_4
XFILLER_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07333_ _07333_/A _07333_/B vssd1 vssd1 vccd1 vccd1 _07333_/X sky130_fd_sc_hd__or2_4
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_118_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10735_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07264_ _07926_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _10400_/D sky130_fd_sc_hd__or2_1
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09003_ _11353_/Q _09013_/B vssd1 vssd1 vccd1 vccd1 _09003_/X sky130_fd_sc_hd__or2_1
X_06215_ _11799_/Q _09154_/A _06697_/B1 _11505_/Q vssd1 vssd1 vccd1 vccd1 _06215_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_118_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07195_ _07211_/A _10358_/Q _07437_/S vssd1 vssd1 vccd1 vccd1 _07195_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06146_ _05704_/X _06665_/A2 _06082_/X _06622_/B2 _06145_/X vssd1 vssd1 vccd1 vccd1
+ _10227_/D sky130_fd_sc_hd__a221o_1
XFILLER_104_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06077_ _06431_/A _06059_/X _06064_/X _06619_/A1 vssd1 vssd1 vccd1 vccd1 _06077_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_67_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout501 _08921_/C1 vssd1 vssd1 vccd1 vccd1 _08947_/C1 sky130_fd_sc_hd__buf_4
Xfanout512 _08816_/A vssd1 vssd1 vccd1 vccd1 _08819_/A sky130_fd_sc_hd__buf_6
X_09905_ _11707_/Q _09565_/B _09950_/B1 _11704_/Q vssd1 vssd1 vccd1 vccd1 _09905_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout523 _07659_/A vssd1 vssd1 vccd1 vccd1 _07476_/A sky130_fd_sc_hd__buf_4
XFILLER_154_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout534 fanout536/X vssd1 vssd1 vccd1 vccd1 _08664_/A sky130_fd_sc_hd__clkbuf_8
Xfanout545 fanout555/X vssd1 vssd1 vccd1 vccd1 _07918_/A sky130_fd_sc_hd__buf_2
Xfanout556 _08773_/A vssd1 vssd1 vccd1 vccd1 _08793_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _11459_/Q _09876_/A2 _09878_/B1 _10780_/Q vssd1 vssd1 vccd1 vccd1 _09836_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout567 _08670_/A vssd1 vssd1 vccd1 vccd1 _08684_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout578 _06898_/Y vssd1 vssd1 vccd1 vccd1 fanout578/X sky130_fd_sc_hd__buf_4
XFILLER_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout589 _06855_/B vssd1 vssd1 vccd1 vccd1 _06535_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06979_ _10257_/Q _06995_/B vssd1 vssd1 vccd1 vccd1 _06979_/X sky130_fd_sc_hd__or2_1
XFILLER_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09767_ _11645_/Q _09766_/X _09770_/S vssd1 vssd1 vccd1 vccd1 _11645_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _11215_/Q _10128_/A0 _08718_/S vssd1 vssd1 vccd1 vccd1 _08719_/B sky130_fd_sc_hd__mux2_1
XFILLER_73_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _11636_/Q _11640_/Q _09702_/S vssd1 vssd1 vccd1 vccd1 _09699_/B sky130_fd_sc_hd__mux2_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _08649_/A _08649_/B _08649_/C vssd1 vssd1 vccd1 vccd1 _08750_/B sky130_fd_sc_hd__and3_4
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _11665_/CLK _11660_/D vssd1 vssd1 vccd1 vccd1 _11660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10611_ _10932_/CLK _10611_/D vssd1 vssd1 vccd1 vccd1 _10611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11591_ _11604_/CLK _11591_/D vssd1 vssd1 vccd1 vccd1 _11591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10542_ _10666_/CLK _10542_/D vssd1 vssd1 vccd1 vccd1 _10542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10473_ _11641_/CLK _10473_/D vssd1 vssd1 vccd1 vccd1 _10473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_4__f_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_4__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11025_ _11186_/CLK _11025_/D vssd1 vssd1 vccd1 vccd1 _11025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10809_ _11473_/CLK _10809_/D vssd1 vssd1 vccd1 vccd1 _10809_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_19 _06431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _11791_/CLK _11789_/D vssd1 vssd1 vccd1 vccd1 _11789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06000_ _06431_/A _06000_/B _06000_/C vssd1 vssd1 vccd1 vccd1 _06000_/X sky130_fd_sc_hd__or3_2
XFILLER_12_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput126 _05716_/X vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_4
Xoutput137 _11617_/Q vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__buf_4
XFILLER_114_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput148 _11571_/Q vssd1 vssd1 vccd1 vccd1 ram_addr[2] sky130_fd_sc_hd__buf_4
Xoutput159 _11579_/Q vssd1 vssd1 vccd1 vccd1 rom_addr[1] sky130_fd_sc_hd__buf_4
XFILLER_130_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07951_ _10793_/Q _07941_/Y _07944_/Y _07333_/X vssd1 vssd1 vccd1 vccd1 _10793_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06902_ _08286_/A _08649_/B _10158_/B vssd1 vssd1 vccd1 vccd1 _06922_/B sky130_fd_sc_hd__and3_4
XFILLER_96_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07882_ _07028_/A _07966_/S _07881_/X _07882_/C1 vssd1 vssd1 vccd1 vccd1 _10759_/D
+ sky130_fd_sc_hd__o211a_1
X_06833_ _11447_/Q _07777_/A _06727_/B _10414_/Q vssd1 vssd1 vccd1 vccd1 _06833_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09621_ _10730_/Q _09567_/B _09570_/B _10799_/Q vssd1 vssd1 vccd1 vccd1 _09621_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09552_ _09552_/A1 _09541_/Y _09551_/X _09447_/B vssd1 vssd1 vccd1 vccd1 _11628_/D
+ sky130_fd_sc_hd__o211a_1
X_06764_ _10763_/Q _07854_/A _06875_/B1 _10674_/Q vssd1 vssd1 vccd1 vccd1 _06764_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_97_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08503_ _11102_/Q _08503_/B vssd1 vssd1 vccd1 vccd1 _08503_/X sky130_fd_sc_hd__or2_1
X_05715_ _11039_/Q _05537_/Y _05573_/Y _11042_/Q _05712_/X vssd1 vssd1 vccd1 vccd1
+ _05716_/D sky130_fd_sc_hd__a221o_2
XFILLER_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ _09515_/B _09515_/C vssd1 vssd1 vccd1 vccd1 _09522_/C sky130_fd_sc_hd__nand2b_1
X_06695_ _06689_/X _06694_/X _06743_/B vssd1 vssd1 vccd1 vccd1 _06695_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08434_ _11059_/Q _08425_/Y _08426_/Y _07095_/X vssd1 vssd1 vccd1 vccd1 _11059_/D
+ sky130_fd_sc_hd__o22a_1
X_05646_ _11290_/Q _05609_/Y _05627_/Y _11285_/Q vssd1 vssd1 vccd1 vccd1 _05655_/A
+ sky130_fd_sc_hd__a22o_1
X_08365_ _09016_/A _08665_/C _10087_/C vssd1 vssd1 vccd1 vccd1 _08365_/X sky130_fd_sc_hd__or3_2
X_05577_ _05631_/A2 _11368_/Q _11364_/Q _05631_/B1 _05575_/X vssd1 vssd1 vccd1 vccd1
+ _05577_/X sky130_fd_sc_hd__a221o_1
X_07316_ _07617_/A _07316_/B vssd1 vssd1 vccd1 vccd1 _07316_/X sky130_fd_sc_hd__or2_4
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08296_ _10982_/Q _07232_/X _08298_/S vssd1 vssd1 vccd1 vccd1 _10982_/D sky130_fd_sc_hd__mux2_1
X_07247_ _07034_/X _07663_/S _07246_/S _10392_/Q _07309_/A vssd1 vssd1 vccd1 vccd1
+ _10392_/D sky130_fd_sc_hd__a221o_1
XFILLER_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07178_ _10350_/Q _09228_/B vssd1 vssd1 vccd1 vccd1 _07178_/X sky130_fd_sc_hd__or2_1
XFILLER_156_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06129_ _10914_/Q _08166_/A _05865_/B _11771_/Q vssd1 vssd1 vccd1 vccd1 _06129_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_156_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_wb_clk_i clkbuf_leaf_88_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11812_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout320 _07259_/S vssd1 vssd1 vccd1 vccd1 _09187_/S sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_15_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11308_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout331 _09240_/S vssd1 vssd1 vccd1 vccd1 _07172_/S sky130_fd_sc_hd__buf_8
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout342 _08243_/X vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__buf_6
Xfanout353 _07022_/X vssd1 vssd1 vccd1 vccd1 _09232_/B2 sky130_fd_sc_hd__buf_12
XFILLER_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout364 _07057_/X vssd1 vssd1 vccd1 vccd1 _07098_/B sky130_fd_sc_hd__buf_6
XFILLER_87_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout375 _08322_/A vssd1 vssd1 vccd1 vccd1 _07309_/A sky130_fd_sc_hd__buf_6
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout386 _07614_/A vssd1 vssd1 vccd1 vccd1 _09193_/A sky130_fd_sc_hd__buf_6
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout397 _07225_/A vssd1 vssd1 vccd1 vccd1 _07005_/A sky130_fd_sc_hd__clkbuf_16
X_09819_ _09825_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _11653_/D sky130_fd_sc_hd__and2_1
XFILLER_98_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11712_/CLK _11712_/D vssd1 vssd1 vccd1 vccd1 _11712_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11661_/CLK _11643_/D vssd1 vssd1 vccd1 vccd1 _11643_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11574_ _11575_/CLK _11574_/D vssd1 vssd1 vccd1 vccd1 _11574_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_126_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput17 rom_value[16] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
Xinput28 rom_value[26] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10525_ _10725_/CLK _10525_/D vssd1 vssd1 vccd1 vccd1 _10525_/Q sky130_fd_sc_hd__dfxtp_1
Xinput39 rom_value[7] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10456_ _11224_/CLK _10456_/D vssd1 vssd1 vccd1 vccd1 _10456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10387_ _11743_/CLK _10387_/D vssd1 vssd1 vccd1 vccd1 _10387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11008_ _11235_/CLK _11008_/D vssd1 vssd1 vccd1 vccd1 _11008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05500_ _10245_/Q input57/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05500_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06480_ _10289_/Q _09325_/A _09248_/A _10320_/Q vssd1 vssd1 vccd1 vccd1 _06480_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05431_ _11151_/Q _11150_/Q _09430_/B vssd1 vssd1 vccd1 vccd1 _05433_/C sky130_fd_sc_hd__mux2_1
XFILLER_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08150_ _10901_/Q _08164_/B vssd1 vssd1 vccd1 vccd1 _08150_/X sky130_fd_sc_hd__or2_1
X_05362_ _05362_/A _05362_/B _05362_/C _05362_/D vssd1 vssd1 vccd1 vccd1 _05368_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07101_ _10306_/Q _07100_/X _07109_/S vssd1 vssd1 vccd1 vccd1 _10306_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08081_ _10866_/Q _08085_/B vssd1 vssd1 vccd1 vccd1 _08081_/X sky130_fd_sc_hd__or2_1
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05293_ _11130_/Q _11129_/Q _05392_/S vssd1 vssd1 vccd1 vccd1 _05296_/B sky130_fd_sc_hd__mux2_1
X_07032_ _10275_/Q _07477_/S _07038_/S _07243_/B vssd1 vssd1 vccd1 vccd1 _07033_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_114_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ _09283_/A1 _08989_/B _09290_/B1 vssd1 vssd1 vccd1 vccd1 _08983_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07934_ _07934_/A _07934_/B vssd1 vssd1 vccd1 vccd1 _10784_/D sky130_fd_sc_hd__or2_1
XFILLER_151_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07865_ _10751_/Q _07883_/B vssd1 vssd1 vccd1 vccd1 _07865_/X sky130_fd_sc_hd__or2_1
XFILLER_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09604_ _10382_/Q _09568_/B _09571_/C _10393_/Q vssd1 vssd1 vccd1 vccd1 _09604_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06816_ _10786_/Q _06875_/A2 _06877_/B1 _10579_/Q _06815_/X vssd1 vssd1 vccd1 vccd1
+ _06816_/X sky130_fd_sc_hd__o221a_1
XFILLER_44_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07796_ _07796_/A _07796_/B vssd1 vssd1 vccd1 vccd1 _10705_/D sky130_fd_sc_hd__or2_1
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06747_ _10490_/Q _06803_/A2 _06856_/A2 _10329_/Q _06746_/X vssd1 vssd1 vccd1 vccd1
+ _06747_/X sky130_fd_sc_hd__o221a_1
XFILLER_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09535_ _09528_/A _09502_/B _09512_/Y _09534_/X _09529_/A vssd1 vssd1 vccd1 vccd1
+ _11622_/D sky130_fd_sc_hd__o311a_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_133_wb_clk_i clkbuf_4_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11710_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09466_ _09475_/A _09464_/X _09465_/Y _09414_/S vssd1 vssd1 vccd1 vccd1 _11599_/D
+ sky130_fd_sc_hd__a22o_1
X_06678_ _11049_/Q _06735_/A2 _06737_/B1 _10971_/Q vssd1 vssd1 vccd1 vccd1 _06678_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05629_ _11790_/Q _05629_/A2 _05629_/B1 _11784_/Q vssd1 vssd1 vccd1 vccd1 _05629_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08417_ _09216_/A0 _08404_/S _08416_/X _08921_/C1 vssd1 vssd1 vccd1 vccd1 _11049_/D
+ sky130_fd_sc_hd__o211a_1
X_09397_ _09971_/A0 _11563_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _11563_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08348_ _09323_/A0 _11017_/Q _08354_/S vssd1 vssd1 vccd1 vccd1 _08349_/B sky130_fd_sc_hd__mux2_1
XFILLER_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08279_ _09216_/A0 _08276_/S _08278_/X _08921_/C1 vssd1 vssd1 vccd1 vccd1 _10971_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10310_ _10727_/CLK _10310_/D vssd1 vssd1 vccd1 vccd1 _10310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11290_ _11291_/CLK _11290_/D vssd1 vssd1 vccd1 vccd1 _11290_/Q sky130_fd_sc_hd__dfxtp_1
X_10241_ _11622_/CLK _10241_/D vssd1 vssd1 vccd1 vccd1 _10241_/Q sky130_fd_sc_hd__dfxtp_2
X_10172_ _10172_/A1 _10176_/B _10178_/B1 vssd1 vssd1 vccd1 vccd1 _10172_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11626_ _11657_/CLK _11626_/D vssd1 vssd1 vccd1 vccd1 _11626_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_129_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11557_ _11675_/CLK _11557_/D vssd1 vssd1 vccd1 vccd1 _11557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10508_ _11665_/CLK _10508_/D vssd1 vssd1 vccd1 vccd1 _10508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11488_ _11497_/CLK _11488_/D vssd1 vssd1 vccd1 vccd1 _11488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10439_ _11177_/CLK _10439_/D vssd1 vssd1 vccd1 vccd1 _10439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05980_ _10282_/Q _07046_/A _06856_/A2 _10313_/Q vssd1 vssd1 vccd1 vccd1 _05980_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07650_ _10614_/Q _07100_/X _07651_/S vssd1 vssd1 vccd1 vccd1 _10614_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06601_ _07083_/A _06601_/B _06601_/C vssd1 vssd1 vccd1 vccd1 _06601_/X sky130_fd_sc_hd__or3_4
XFILLER_66_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07581_ _07932_/A1 _10574_/Q _07593_/S vssd1 vssd1 vccd1 vccd1 _07582_/B sky130_fd_sc_hd__mux2_1
X_09320_ _10114_/A0 _11513_/Q _09324_/S vssd1 vssd1 vccd1 vccd1 _11513_/D sky130_fd_sc_hd__mux2_1
X_06532_ _11164_/Q _06649_/A2 _06528_/X _06531_/X vssd1 vssd1 vccd1 vccd1 _06532_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_59_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09251_ _10088_/A1 _09249_/X _09250_/X _10155_/C1 vssd1 vssd1 vccd1 vccd1 _11478_/D
+ sky130_fd_sc_hd__o211a_1
X_06463_ _10448_/Q _06635_/A2 _08647_/B _10307_/Q vssd1 vssd1 vccd1 vccd1 _06467_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_61_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08202_ _08839_/A _08202_/B vssd1 vssd1 vccd1 vccd1 _10935_/D sky130_fd_sc_hd__or2_1
XFILLER_138_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05414_ _10422_/Q _10421_/Q _05414_/S vssd1 vssd1 vccd1 vccd1 _05417_/B sky130_fd_sc_hd__mux2_1
X_09182_ _09182_/A0 _11436_/Q _09184_/S vssd1 vssd1 vccd1 vccd1 _09182_/X sky130_fd_sc_hd__mux2_1
X_06394_ _10817_/Q _06639_/B1 _06640_/B1 _11140_/Q vssd1 vssd1 vccd1 vccd1 _06394_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08133_ _08835_/A _08133_/B vssd1 vssd1 vccd1 vccd1 _10892_/D sky130_fd_sc_hd__or2_1
XFILLER_105_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05345_ _05345_/A _05345_/B _05345_/C _05345_/D vssd1 vssd1 vccd1 vccd1 _05346_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_147_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08064_ _08835_/A _08064_/B vssd1 vssd1 vccd1 vccd1 _10857_/D sky130_fd_sc_hd__or2_1
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05276_ _10452_/Q _10451_/Q _05391_/S vssd1 vssd1 vccd1 vccd1 _05280_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07015_ _07015_/A _07107_/B vssd1 vssd1 vccd1 vccd1 _07095_/B sky130_fd_sc_hd__and2_4
XFILLER_66_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08966_ _11334_/Q _08965_/A _08965_/Y _09833_/A vssd1 vssd1 vccd1 vccd1 _11334_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07917_ _08846_/A0 _10776_/Q _09218_/S vssd1 vssd1 vccd1 vccd1 _07918_/B sky130_fd_sc_hd__mux2_1
XFILLER_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08897_ _11306_/Q _07013_/X _08901_/S vssd1 vssd1 vccd1 vccd1 _11306_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07848_ _08810_/A _08726_/S vssd1 vssd1 vccd1 vccd1 _07852_/S sky130_fd_sc_hd__nor2_8
XFILLER_29_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07779_ _07303_/A _10697_/Q _07817_/S vssd1 vssd1 vccd1 vccd1 _07780_/B sky130_fd_sc_hd__mux2_1
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09518_ _09492_/B _09528_/B _09516_/Y _09517_/X _09825_/A vssd1 vssd1 vccd1 vccd1
+ _11615_/D sky130_fd_sc_hd__o311a_1
X_10790_ _11234_/CLK _10790_/D vssd1 vssd1 vccd1 vccd1 _10790_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09441_/B input19/X _09441_/A vssd1 vssd1 vccd1 vccd1 _09449_/X sky130_fd_sc_hd__o21a_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _11411_/CLK _11411_/D vssd1 vssd1 vccd1 vccd1 _11411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11342_ _11495_/CLK _11342_/D vssd1 vssd1 vccd1 vccd1 _11342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11023_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11273_ _11634_/CLK _11273_/D vssd1 vssd1 vccd1 vccd1 _11273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10224_ _10644_/CLK _10224_/D vssd1 vssd1 vccd1 vccd1 _10224_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10155_ _10177_/A1 _10137_/X _10154_/X _10155_/C1 vssd1 vssd1 vccd1 vccd1 _11790_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10086_ _10086_/A _10158_/B _10136_/C vssd1 vssd1 vccd1 vccd1 _10104_/B sky130_fd_sc_hd__and3_4
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10988_ _11633_/CLK _10988_/D vssd1 vssd1 vccd1 vccd1 _10988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11609_ _11663_/CLK _11609_/D vssd1 vssd1 vccd1 vccd1 _11609_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05130_ _10611_/Q _10610_/Q _05391_/S vssd1 vssd1 vccd1 vccd1 _05134_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout908 _06852_/A1 vssd1 vssd1 vccd1 vccd1 _06853_/A1 sky130_fd_sc_hd__buf_4
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout919 _06651_/C1 vssd1 vssd1 vccd1 vccd1 _06808_/C1 sky130_fd_sc_hd__buf_6
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _11268_/Q _10135_/A0 _08820_/S vssd1 vssd1 vccd1 vccd1 _08821_/B sky130_fd_sc_hd__mux2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05963_ _11669_/Q _09965_/A _08311_/A _10994_/Q vssd1 vssd1 vccd1 vccd1 _05963_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08751_ _08469_/A _08748_/S _08750_/X _08578_/A vssd1 vssd1 vccd1 vccd1 _11232_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07702_ _10650_/Q _07693_/Y _07697_/Y _09232_/B2 vssd1 vssd1 vccd1 vccd1 _10650_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05894_ _11391_/Q _09082_/A _09110_/A _11404_/Q vssd1 vssd1 vccd1 vccd1 _05894_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_113_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08682_ _08682_/A _08682_/B vssd1 vssd1 vccd1 vccd1 _11195_/D sky130_fd_sc_hd__or2_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07633_ _10602_/Q _08326_/B2 _07637_/S vssd1 vssd1 vccd1 vccd1 _10602_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07564_ _07916_/A _07564_/B vssd1 vssd1 vccd1 vccd1 _10565_/D sky130_fd_sc_hd__or2_1
XFILLER_59_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09303_ _11502_/Q _09293_/X _09302_/X vssd1 vssd1 vccd1 vccd1 _11502_/D sky130_fd_sc_hd__a21o_1
X_06515_ _06512_/X _06514_/X _07083_/A vssd1 vssd1 vccd1 vccd1 _06515_/X sky130_fd_sc_hd__a21o_2
XFILLER_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07495_ _07451_/X _10531_/Q _07496_/S vssd1 vssd1 vccd1 vccd1 _10531_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09234_ _09234_/A0 _11468_/Q _09243_/C vssd1 vssd1 vccd1 vccd1 _09234_/X sky130_fd_sc_hd__mux2_1
X_06446_ _11113_/Q _06646_/A2 _06444_/X _06445_/X vssd1 vssd1 vccd1 vccd1 _06446_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09165_ _11427_/Q _09171_/B vssd1 vssd1 vccd1 vccd1 _09165_/X sky130_fd_sc_hd__or2_1
X_06377_ _11161_/Q _06735_/B1 _06737_/B1 _10964_/Q vssd1 vssd1 vccd1 vccd1 _06377_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08116_ _08193_/A _08116_/B vssd1 vssd1 vccd1 vccd1 _10884_/D sky130_fd_sc_hd__or2_1
XFILLER_107_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05328_ _10460_/Q _10459_/Q _05382_/S vssd1 vssd1 vccd1 vccd1 _05329_/D sky130_fd_sc_hd__mux2_1
X_09096_ _09285_/A1 _09082_/X _09095_/X _09279_/C1 vssd1 vssd1 vccd1 vccd1 _11395_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08047_ _08749_/A _08047_/B vssd1 vssd1 vccd1 vccd1 _10849_/D sky130_fd_sc_hd__or2_1
X_05259_ _05259_/A _05259_/B vssd1 vssd1 vccd1 vccd1 _05259_/Y sky130_fd_sc_hd__nor2_8
XFILLER_153_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09998_ _09998_/A _10108_/B _10119_/C vssd1 vssd1 vccd1 vccd1 _10008_/S sky130_fd_sc_hd__or3_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08949_ _09668_/B _09488_/C _09668_/D vssd1 vssd1 vccd1 vccd1 _08958_/A sky130_fd_sc_hd__nor3_2
XFILLER_69_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _11766_/CLK _10911_/D vssd1 vssd1 vccd1 vccd1 _10911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10842_ _11527_/CLK _10842_/D vssd1 vssd1 vccd1 vccd1 _10842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10773_ _10773_/CLK _10773_/D vssd1 vssd1 vccd1 vccd1 _10773_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11325_ _11325_/CLK _11325_/D vssd1 vssd1 vccd1 vccd1 _11325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11256_ _11812_/CLK _11256_/D vssd1 vssd1 vccd1 vccd1 _11256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _11808_/CLK _10207_/D vssd1 vssd1 vccd1 vccd1 _10207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11187_ _11607_/CLK _11187_/D vssd1 vssd1 vccd1 vccd1 _11187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10138_ _11782_/Q _10154_/B vssd1 vssd1 vccd1 vccd1 _10138_/X sky130_fd_sc_hd__or2_1
XFILLER_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10069_ _10080_/A0 _11730_/Q _10071_/S vssd1 vssd1 vccd1 vccd1 _11730_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06300_ _10661_/Q _07455_/A vssd1 vssd1 vccd1 vccd1 _06300_/X sky130_fd_sc_hd__or2_1
XFILLER_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07280_ _07926_/A _07280_/B vssd1 vssd1 vccd1 vccd1 _10408_/D sky130_fd_sc_hd__or2_1
XFILLER_143_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06231_ _11809_/Q _10180_/A _06229_/X _06230_/X vssd1 vssd1 vccd1 vccd1 _06231_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06162_ _11093_/Q _08472_/A _06158_/X _06161_/X vssd1 vssd1 vccd1 vccd1 _06162_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05113_ _05113_/A _05113_/B vssd1 vssd1 vccd1 vccd1 _05113_/Y sky130_fd_sc_hd__nor2_8
XFILLER_89_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06093_ _07297_/A _06093_/B _06093_/C vssd1 vssd1 vccd1 vccd1 _06093_/X sky130_fd_sc_hd__or3_2
XFILLER_132_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09921_ _10478_/Q _09568_/B _09566_/B _10476_/Q vssd1 vssd1 vccd1 vccd1 _09921_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout705 _11587_/Q vssd1 vssd1 vccd1 vccd1 _09540_/A sky130_fd_sc_hd__buf_12
Xfanout716 fanout726/X vssd1 vssd1 vccd1 vccd1 _06556_/B1 sky130_fd_sc_hd__buf_4
Xfanout727 _06871_/B1 vssd1 vssd1 vccd1 vccd1 _06710_/B sky130_fd_sc_hd__buf_6
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _11449_/Q _09909_/A2 _09565_/C _10708_/Q vssd1 vssd1 vccd1 vccd1 _09852_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout738 _05751_/X vssd1 vssd1 vccd1 vccd1 fanout738/X sky130_fd_sc_hd__buf_12
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 fanout755/X vssd1 vssd1 vccd1 vccd1 _08472_/A sky130_fd_sc_hd__buf_4
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08803_ _08869_/A _08803_/B vssd1 vssd1 vccd1 vccd1 _11257_/D sky130_fd_sc_hd__or2_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _05372_/S _09672_/B _09674_/A _11590_/Q vssd1 vssd1 vccd1 vccd1 _09783_/X
+ sky130_fd_sc_hd__o22a_1
X_06995_ _10265_/Q _06995_/B vssd1 vssd1 vccd1 vccd1 _06995_/X sky130_fd_sc_hd__or2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08734_ _11224_/Q _08750_/B vssd1 vssd1 vccd1 vccd1 _08734_/X sky130_fd_sc_hd__or2_1
XFILLER_113_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05946_ _06633_/A _05939_/X _05944_/X _06619_/A1 _05934_/X vssd1 vssd1 vccd1 vccd1
+ _05946_/X sky130_fd_sc_hd__o311a_1
XFILLER_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08665_ _08665_/A _09249_/A _08665_/C _10087_/C vssd1 vssd1 vccd1 vccd1 _08665_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_22_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_109 fanout793/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05877_ _11054_/Q _08054_/A _08123_/A _11172_/Q _06392_/C1 vssd1 vssd1 vccd1 vccd1
+ _05877_/X sky130_fd_sc_hd__o221a_1
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _10592_/Q _07613_/Y _07614_/Y _07227_/X vssd1 vssd1 vccd1 vccd1 _10592_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08596_ _08873_/A _08596_/B vssd1 vssd1 vccd1 vccd1 _11152_/D sky130_fd_sc_hd__or2_1
XFILLER_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07547_ _07785_/A0 _10557_/Q _07591_/S vssd1 vssd1 vccd1 vccd1 _07548_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07478_ _10043_/A _07478_/B vssd1 vssd1 vccd1 vccd1 _10517_/D sky130_fd_sc_hd__or2_1
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09217_ _07922_/A _09216_/X _09243_/B vssd1 vssd1 vccd1 vccd1 _11457_/D sky130_fd_sc_hd__o21a_1
X_06429_ _10618_/Q _06642_/A2 _06428_/X _06642_/C1 vssd1 vssd1 vccd1 vccd1 _06429_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09148_ _11419_/Q _09132_/X _09147_/X vssd1 vssd1 vccd1 vccd1 _11419_/D sky130_fd_sc_hd__a21o_1
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09079_ _10178_/A1 _09077_/B _08783_/A vssd1 vssd1 vccd1 vccd1 _09079_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11110_ _11329_/CLK _11110_/D vssd1 vssd1 vccd1 vccd1 _11110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_3__f_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_3__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11041_ _11243_/CLK _11041_/D vssd1 vssd1 vccd1 vccd1 _11041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ input75/X vssd1 vssd1 vccd1 vccd1 _11874_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ _11634_/CLK _10825_/D vssd1 vssd1 vccd1 vccd1 _10825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10756_ _10782_/CLK _10756_/D vssd1 vssd1 vccd1 vccd1 _10756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ _11661_/CLK _10687_/D vssd1 vssd1 vccd1 vccd1 _10687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11308_ _11308_/CLK _11308_/D vssd1 vssd1 vccd1 vccd1 _11308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11239_ _11411_/CLK _11239_/D vssd1 vssd1 vccd1 vccd1 _11239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05800_ _10607_/Q _06468_/B _06152_/B _10610_/Q _07083_/B vssd1 vssd1 vccd1 vccd1
+ _05800_/X sky130_fd_sc_hd__o221a_2
X_06780_ _10784_/Q _06875_/A2 _06779_/X _06878_/C1 vssd1 vssd1 vccd1 vccd1 _06780_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05731_ _06450_/A _10222_/Q vssd1 vssd1 vccd1 vccd1 _05731_/X sky130_fd_sc_hd__and2_1
XFILLER_76_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05662_ _11244_/Q _05609_/Y _05627_/Y _11239_/Q vssd1 vssd1 vccd1 vccd1 _05662_/X
+ sky130_fd_sc_hd__a22o_1
X_08450_ _11071_/Q _07623_/X _07628_/S _07090_/A vssd1 vssd1 vccd1 vccd1 _11071_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07401_ _07010_/A _10477_/Q _07429_/S vssd1 vssd1 vccd1 vccd1 _07402_/B sky130_fd_sc_hd__mux2_1
X_08381_ _08665_/A _08365_/X _08380_/Y _09032_/C1 vssd1 vssd1 vccd1 vccd1 _11032_/D
+ sky130_fd_sc_hd__o211a_1
X_05593_ _05629_/A2 _11486_/Q _11480_/Q _05629_/B1 vssd1 vssd1 vccd1 vccd1 _05593_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07332_ _10432_/Q _07323_/Y _07325_/Y _07318_/X vssd1 vssd1 vccd1 vccd1 _10432_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07263_ _10021_/A0 _10400_/Q _07277_/S vssd1 vssd1 vccd1 vccd1 _07264_/B sky130_fd_sc_hd__mux2_1
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06214_ _11753_/Q _10087_/A _06214_/B1 _11789_/Q _06214_/C1 vssd1 vssd1 vccd1 vccd1
+ _06214_/X sky130_fd_sc_hd__o221a_2
XFILLER_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09002_ _11352_/Q _08994_/X _09001_/X vssd1 vssd1 vccd1 vccd1 _11352_/D sky130_fd_sc_hd__a21o_1
X_07194_ _08661_/A _07429_/S _07192_/Y _10357_/Q _08439_/A vssd1 vssd1 vccd1 vccd1
+ _10357_/D sky130_fd_sc_hd__o221a_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06145_ _06855_/B _06082_/X _06144_/X _05819_/B vssd1 vssd1 vccd1 vccd1 _06145_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06076_ _07151_/B _06049_/X _06054_/X _06039_/X vssd1 vssd1 vccd1 vccd1 _06076_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_63_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09904_ _11705_/Q _09573_/B _09572_/C _11720_/Q _09903_/X vssd1 vssd1 vccd1 vccd1
+ _09907_/C sky130_fd_sc_hd__a221o_1
Xfanout502 _09048_/C1 vssd1 vssd1 vccd1 vccd1 _08921_/C1 sky130_fd_sc_hd__buf_4
Xfanout513 _08196_/A vssd1 vssd1 vccd1 vccd1 _08193_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout524 _07659_/A vssd1 vssd1 vccd1 vccd1 _08733_/A sky130_fd_sc_hd__buf_4
Xfanout535 fanout536/X vssd1 vssd1 vccd1 vccd1 _08757_/A sky130_fd_sc_hd__buf_8
XFILLER_154_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout546 _07922_/A vssd1 vssd1 vccd1 vccd1 _07930_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _10777_/Q _09873_/B1 _09875_/B1 _11452_/Q _09834_/X vssd1 vssd1 vccd1 vccd1
+ _09842_/A sky130_fd_sc_hd__a221o_2
XFILLER_59_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout557 _08773_/A vssd1 vssd1 vccd1 vccd1 _08847_/A sky130_fd_sc_hd__buf_6
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout568 _08670_/A vssd1 vssd1 vccd1 vccd1 _08536_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout579 _05819_/Y vssd1 vssd1 vccd1 vccd1 _06622_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_100_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09766_ input8/X _09740_/Y _09765_/X vssd1 vssd1 vccd1 vccd1 _09766_/X sky130_fd_sc_hd__a21o_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06978_ _10088_/A1 _06976_/X _06977_/X _06990_/C1 vssd1 vssd1 vccd1 vccd1 _10256_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08717_ _11214_/Q _08726_/S _07852_/S _08811_/B2 vssd1 vssd1 vccd1 vccd1 _11214_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05929_ _10437_/Q _06634_/B1 _07111_/A _11768_/Q vssd1 vssd1 vccd1 vccd1 _05929_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09697_ _09703_/A _09697_/B vssd1 vssd1 vccd1 vccd1 _11639_/D sky130_fd_sc_hd__or2_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _11180_/Q _08645_/S _08647_/X _08821_/A vssd1 vssd1 vccd1 vccd1 _11180_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _08579_/A0 _11145_/Q _08589_/S vssd1 vssd1 vccd1 vccd1 _08580_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10610_ _10932_/CLK _10610_/D vssd1 vssd1 vccd1 vccd1 _10610_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11590_ _11652_/CLK _11590_/D vssd1 vssd1 vccd1 vccd1 _11590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ _11472_/CLK _10541_/D vssd1 vssd1 vccd1 vccd1 _10541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10472_ _11641_/CLK _10472_/D vssd1 vssd1 vccd1 vccd1 _10472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11024_ _11733_/CLK _11024_/D vssd1 vssd1 vccd1 vccd1 _11024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10808_ _10808_/CLK _10808_/D vssd1 vssd1 vccd1 vccd1 _10808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11788_ _11791_/CLK _11788_/D vssd1 vssd1 vccd1 vccd1 _11788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10739_ _11766_/CLK _10739_/D vssd1 vssd1 vccd1 vccd1 _10739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput127 _05728_/X vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_4
XFILLER_126_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput138 _11618_/Q vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__buf_4
Xoutput149 _11572_/Q vssd1 vssd1 vccd1 vccd1 ram_addr[3] sky130_fd_sc_hd__buf_4
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07950_ _10792_/Q _07942_/Y _07943_/Y _07314_/X vssd1 vssd1 vccd1 vccd1 _10792_/D
+ sky130_fd_sc_hd__o22a_1
X_06901_ _06901_/A _08243_/C _08243_/D vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__or3_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07881_ _10759_/Q _07893_/B vssd1 vssd1 vccd1 vccd1 _07881_/X sky130_fd_sc_hd__or2_1
XFILLER_60_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09620_ _10796_/Q _09566_/C _09566_/D _10736_/Q vssd1 vssd1 vccd1 vccd1 _09620_/X
+ sky130_fd_sc_hd__a22o_1
X_06832_ _10502_/Q _07440_/A vssd1 vssd1 vccd1 vccd1 _06832_/X sky130_fd_sc_hd__or2_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09551_ _11630_/Q _09538_/X _09542_/X vssd1 vssd1 vccd1 vccd1 _09551_/X sky130_fd_sc_hd__a21o_1
X_06763_ _11458_/Q _06875_/A2 _07254_/A _11437_/Q vssd1 vssd1 vccd1 vccd1 _06763_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08502_ _08757_/A _08502_/B vssd1 vssd1 vccd1 vccd1 _11101_/D sky130_fd_sc_hd__or2_1
XFILLER_3_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05714_ _11048_/Q _05561_/Y _05585_/Y _11047_/Q _05713_/X vssd1 vssd1 vccd1 vccd1
+ _05716_/C sky130_fd_sc_hd__a221o_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06694_ _10500_/Q _06728_/B1 _06690_/X _06693_/X vssd1 vssd1 vccd1 vccd1 _06694_/X
+ sky130_fd_sc_hd__o211a_2
X_09482_ _08951_/X _09481_/Y _09959_/A vssd1 vssd1 vccd1 vccd1 _11604_/D sky130_fd_sc_hd__a21oi_1
XFILLER_51_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08433_ _11058_/Q _08424_/Y _08427_/Y _07617_/X vssd1 vssd1 vccd1 vccd1 _11058_/D
+ sky130_fd_sc_hd__a22o_1
X_05645_ _11300_/Q _05561_/Y _05585_/Y _11299_/Q vssd1 vssd1 vccd1 vccd1 _05645_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05576_ _05630_/A2 _11362_/Q _11359_/Q _05079_/A _05574_/X vssd1 vssd1 vccd1 vccd1
+ _05579_/A sky130_fd_sc_hd__a221o_4
X_08364_ _08649_/A _08649_/C _10136_/C vssd1 vssd1 vccd1 vccd1 _08438_/B sky130_fd_sc_hd__and3_2
XFILLER_108_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07315_ _10424_/Q _07302_/Y _07305_/Y _07314_/X vssd1 vssd1 vccd1 vccd1 _10424_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08295_ _10981_/Q _07016_/X _08298_/S vssd1 vssd1 vccd1 vccd1 _10981_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07246_ _07245_/X _10391_/Q _07246_/S vssd1 vssd1 vccd1 vccd1 _10391_/D sky130_fd_sc_hd__mux2_1
X_07177_ _08423_/A1 _07172_/S _07176_/X _07884_/C1 vssd1 vssd1 vccd1 vccd1 _10349_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06128_ _10440_/Q _06634_/B1 _06731_/B1 _11074_/Q _06550_/C1 vssd1 vssd1 vccd1 vccd1
+ _06128_/X sky130_fd_sc_hd__o221a_1
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06059_ _06059_/A _06059_/B vssd1 vssd1 vccd1 vccd1 _06059_/X sky130_fd_sc_hd__and2_2
Xfanout310 _07752_/B vssd1 vssd1 vccd1 vccd1 _07750_/B sky130_fd_sc_hd__clkbuf_8
Xfanout321 _07259_/S vssd1 vssd1 vccd1 vccd1 _09184_/S sky130_fd_sc_hd__buf_8
Xfanout332 _07150_/A2 vssd1 vssd1 vccd1 vccd1 _07126_/B sky130_fd_sc_hd__buf_6
Xfanout343 _07324_/X vssd1 vssd1 vccd1 vccd1 _08440_/B2 sky130_fd_sc_hd__buf_12
Xfanout354 _07005_/X vssd1 vssd1 vccd1 vccd1 _08326_/B2 sky130_fd_sc_hd__clkbuf_16
XFILLER_115_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout365 _07057_/X vssd1 vssd1 vccd1 vccd1 _07314_/B sky130_fd_sc_hd__clkbuf_8
Xfanout376 _08902_/B vssd1 vssd1 vccd1 vccd1 _08655_/B sky130_fd_sc_hd__buf_6
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout387 _07614_/A vssd1 vssd1 vccd1 vccd1 _09241_/B1 sky130_fd_sc_hd__buf_4
X_09818_ _09515_/C _09817_/Y _09824_/S vssd1 vssd1 vccd1 vccd1 _09819_/B sky130_fd_sc_hd__mux2_1
Xfanout398 _05434_/Y vssd1 vssd1 vccd1 vccd1 _09572_/D sky130_fd_sc_hd__buf_6
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_55_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11234_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09749_ _09749_/A _09749_/B _09749_/C _09749_/D vssd1 vssd1 vccd1 vccd1 _09757_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_62_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11711_/CLK _11711_/D vssd1 vssd1 vccd1 vccd1 _11711_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11652_/CLK _11642_/D vssd1 vssd1 vccd1 vccd1 _11642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11573_ _11573_/CLK _11573_/D vssd1 vssd1 vccd1 vccd1 _11573_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput18 rom_value[17] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput29 rom_value[27] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_2
X_10524_ _10812_/CLK _10524_/D vssd1 vssd1 vccd1 vccd1 _10524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10455_ _11308_/CLK _10455_/D vssd1 vssd1 vccd1 vccd1 _10455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10386_ _11133_/CLK _10386_/D vssd1 vssd1 vccd1 vccd1 _10386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _11234_/CLK _11007_/D vssd1 vssd1 vccd1 vccd1 _11007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05430_ _10653_/Q _10652_/Q _05430_/S vssd1 vssd1 vccd1 vccd1 _05433_/B sky130_fd_sc_hd__mux2_1
XFILLER_33_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05361_ _11270_/Q _11269_/Q _05372_/S vssd1 vssd1 vccd1 vccd1 _05362_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07100_ _07318_/A _07316_/B vssd1 vssd1 vccd1 vccd1 _07100_/X sky130_fd_sc_hd__or2_4
XFILLER_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08080_ _08761_/A _08080_/B vssd1 vssd1 vccd1 vccd1 _10865_/D sky130_fd_sc_hd__or2_1
X_05292_ _10448_/Q _11132_/Q _05385_/S vssd1 vssd1 vccd1 vccd1 _05296_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07031_ _07031_/A _07928_/A vssd1 vssd1 vccd1 vccd1 _07243_/B sky130_fd_sc_hd__or2_4
X_08982_ _09280_/A1 _08972_/X _08981_/X _09279_/C1 vssd1 vssd1 vccd1 vccd1 _11343_/D
+ sky130_fd_sc_hd__o211a_1
X_07933_ _07933_/A0 _10784_/Q _09221_/C vssd1 vssd1 vccd1 vccd1 _07934_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07864_ _10017_/A0 _07871_/S _07863_/X _07866_/C1 vssd1 vssd1 vccd1 vccd1 _10750_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09603_ _10381_/Q _09566_/C _09566_/D _10630_/Q vssd1 vssd1 vccd1 vccd1 _09603_/X
+ sky130_fd_sc_hd__a22o_1
X_06815_ _10809_/Q _07854_/A _06875_/B1 _10678_/Q vssd1 vssd1 vccd1 vccd1 _06815_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07795_ _08876_/A0 _10705_/Q _07817_/S vssd1 vssd1 vccd1 vccd1 _07796_/B sky130_fd_sc_hd__mux2_1
X_09534_ _09492_/B _09500_/B _09512_/A _11622_/Q vssd1 vssd1 vccd1 vccd1 _09534_/X
+ sky130_fd_sc_hd__a31o_1
X_06746_ _10295_/Q _06873_/A2 _06685_/B _11715_/Q _06745_/X vssd1 vssd1 vccd1 vccd1
+ _06746_/X sky130_fd_sc_hd__o221a_1
XFILLER_97_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09465_ _09679_/B _09478_/A vssd1 vssd1 vccd1 vccd1 _09465_/Y sky130_fd_sc_hd__nand2_1
X_06677_ _11205_/Q _06736_/A2 _08765_/A _11255_/Q vssd1 vssd1 vccd1 vccd1 _06677_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08416_ _11049_/Q _08422_/B vssd1 vssd1 vccd1 vccd1 _08416_/X sky130_fd_sc_hd__or2_1
X_05628_ _11789_/Q _05628_/A2 _05628_/B1 _11786_/Q vssd1 vssd1 vccd1 vccd1 _05628_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09396_ _09396_/A0 _11562_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _11562_/D sky130_fd_sc_hd__mux2_1
XFILLER_123_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08347_ _08492_/A _08347_/B vssd1 vssd1 vccd1 vccd1 _11016_/D sky130_fd_sc_hd__or2_1
XFILLER_138_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05559_ _05619_/A1 _11348_/Q _11344_/Q _05619_/B2 _05557_/X vssd1 vssd1 vccd1 vccd1
+ _05559_/X sky130_fd_sc_hd__a221o_1
XFILLER_123_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _10773_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08278_ _10971_/Q _08284_/B vssd1 vssd1 vccd1 vccd1 _08278_/X sky130_fd_sc_hd__or2_1
X_07229_ _07617_/A _07229_/B vssd1 vssd1 vccd1 vccd1 _07229_/X sky130_fd_sc_hd__or2_4
XFILLER_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10240_ _11663_/CLK _10240_/D vssd1 vssd1 vccd1 vccd1 _10240_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10171_ _10171_/A1 _10159_/X _10170_/X _10177_/C1 vssd1 vssd1 vccd1 vccd1 _11797_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _11657_/CLK _11625_/D vssd1 vssd1 vccd1 vccd1 _11625_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11556_ _11758_/CLK _11556_/D vssd1 vssd1 vccd1 vccd1 _11556_/Q sky130_fd_sc_hd__dfxtp_1
X_10507_ _11743_/CLK _10507_/D vssd1 vssd1 vccd1 vccd1 _10507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11487_ _11809_/CLK _11487_/D vssd1 vssd1 vccd1 vccd1 _11487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10438_ _11268_/CLK _10438_/D vssd1 vssd1 vccd1 vccd1 _10438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _11713_/CLK _10369_/D vssd1 vssd1 vccd1 vccd1 _10369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06600_ _10851_/Q _06643_/A2 _06596_/X _06599_/X vssd1 vssd1 vccd1 vccd1 _06601_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07580_ _07922_/A _07580_/B vssd1 vssd1 vccd1 vccd1 _10573_/D sky130_fd_sc_hd__or2_1
XFILLER_53_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06531_ _11115_/Q _06646_/A2 _06529_/X _06530_/X vssd1 vssd1 vccd1 vccd1 _06531_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_34_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11220_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09250_ _11478_/Q _09266_/B vssd1 vssd1 vccd1 vccd1 _09250_/X sky130_fd_sc_hd__or2_1
XFILLER_34_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06462_ _06453_/X _06454_/X _06456_/X _06633_/A vssd1 vssd1 vccd1 vccd1 _06462_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08201_ _09999_/A0 _10935_/Q _08225_/S vssd1 vssd1 vccd1 vccd1 _08202_/B sky130_fd_sc_hd__mux2_1
X_05413_ _10426_/Q _10425_/Q _05413_/S vssd1 vssd1 vccd1 vccd1 _05417_/A sky130_fd_sc_hd__mux2_1
X_06393_ _10882_/Q _06468_/B _06152_/B _10930_/Q vssd1 vssd1 vccd1 vccd1 _06393_/X
+ sky130_fd_sc_hd__o22a_1
X_09181_ _11435_/Q _09175_/Y _09176_/Y _07333_/X vssd1 vssd1 vccd1 vccd1 _11435_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08132_ _09971_/A0 _10892_/Q _08146_/S vssd1 vssd1 vccd1 vccd1 _08133_/B sky130_fd_sc_hd__mux2_1
X_05344_ _11096_/Q _11095_/Q _05432_/S vssd1 vssd1 vccd1 vccd1 _05345_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05275_ _05275_/A _05275_/B _05275_/C _05275_/D vssd1 vssd1 vccd1 vccd1 _05281_/A
+ sky130_fd_sc_hd__or4_4
X_08063_ _08834_/A0 _10857_/Q _08427_/B vssd1 vssd1 vccd1 vccd1 _08064_/B sky130_fd_sc_hd__mux2_1
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07014_ _10268_/Q _07013_/X _07038_/S vssd1 vssd1 vccd1 vccd1 _10268_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_1335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08965_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _08965_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07916_ _07916_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _10775_/D sky130_fd_sc_hd__or2_1
XFILLER_97_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08896_ _11305_/Q _07008_/X _08901_/S vssd1 vssd1 vccd1 vccd1 _11305_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07847_ _08560_/A _08560_/C _07847_/C vssd1 vssd1 vccd1 vccd1 _08718_/S sky130_fd_sc_hd__and3_4
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07778_ _07778_/A _07854_/B vssd1 vssd1 vccd1 vccd1 _07778_/X sky130_fd_sc_hd__or2_1
XFILLER_44_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09517_ _09525_/A _09489_/C _09516_/A _11615_/Q vssd1 vssd1 vccd1 vccd1 _09517_/X
+ sky130_fd_sc_hd__a31o_1
X_06729_ _10761_/Q _07854_/A _06875_/B1 _10672_/Q _06727_/X vssd1 vssd1 vccd1 vccd1
+ _06729_/X sky130_fd_sc_hd__o221a_1
XFILLER_71_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _09407_/B _09446_/X _09447_/Y _09414_/S vssd1 vssd1 vccd1 vccd1 _11595_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09379_ _11547_/Q _09359_/X _09378_/X vssd1 vssd1 vccd1 vccd1 _11547_/D sky130_fd_sc_hd__a21o_1
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ _11410_/CLK _11410_/D vssd1 vssd1 vccd1 vccd1 _11410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11341_ _11497_/CLK _11341_/D vssd1 vssd1 vccd1 vccd1 _11341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11272_ _11601_/CLK _11272_/D vssd1 vssd1 vccd1 vccd1 _11272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10223_ _10644_/CLK _10223_/D vssd1 vssd1 vccd1 vccd1 _10223_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11385_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10154_ _11790_/Q _10154_/B vssd1 vssd1 vccd1 vccd1 _10154_/X sky130_fd_sc_hd__or2_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10085_ _11745_/Q _07043_/X _10085_/S vssd1 vssd1 vccd1 vccd1 _11745_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10987_ _11633_/CLK _10987_/D vssd1 vssd1 vccd1 vccd1 _10987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11608_ _11811_/CLK _11608_/D vssd1 vssd1 vccd1 vccd1 _11608_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11539_ _11800_/CLK _11539_/D vssd1 vssd1 vccd1 vccd1 _11539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout909 _06577_/A vssd1 vssd1 vccd1 vccd1 _06852_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _11232_/Q _08750_/B vssd1 vssd1 vccd1 vccd1 _08750_/X sky130_fd_sc_hd__or2_1
XFILLER_85_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05962_ _07297_/A _05962_/B _05962_/C vssd1 vssd1 vccd1 vccd1 _05962_/X sky130_fd_sc_hd__or3_4
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07701_ _10649_/Q _07694_/Y _07696_/Y _07232_/X vssd1 vssd1 vccd1 vccd1 _10649_/D
+ sky130_fd_sc_hd__o22a_1
X_08681_ _09124_/A1 _11195_/Q _08707_/S vssd1 vssd1 vccd1 vccd1 _08682_/B sky130_fd_sc_hd__mux2_1
X_05893_ _11490_/Q _08907_/A _08855_/A _11414_/Q _06670_/D1 vssd1 vssd1 vccd1 vccd1
+ _05893_/X sky130_fd_sc_hd__o221a_1
XFILLER_96_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07632_ _10601_/Q _07088_/X _07637_/S vssd1 vssd1 vccd1 vccd1 _10601_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07563_ _08931_/A1 _10565_/Q _07593_/S vssd1 vssd1 vccd1 vccd1 _07564_/B sky130_fd_sc_hd__mux2_1
X_09302_ _10168_/A1 _09310_/B _10178_/B1 vssd1 vssd1 vccd1 vccd1 _09302_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06514_ _11265_/Q _06514_/A2 _05865_/B _11778_/Q _06513_/X vssd1 vssd1 vccd1 vccd1
+ _06514_/X sky130_fd_sc_hd__o221a_1
X_07494_ _10530_/Q _07496_/S _07143_/X _07078_/B _07451_/A vssd1 vssd1 vccd1 vccd1
+ _10530_/D sky130_fd_sc_hd__a221o_1
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09233_ _11467_/Q _09227_/Y _09228_/Y _07318_/X vssd1 vssd1 vccd1 vccd1 _11467_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06445_ _11199_/Q _06645_/A2 _09109_/A _11249_/Q vssd1 vssd1 vccd1 vccd1 _06445_/X
+ sky130_fd_sc_hd__a22o_1
X_09164_ _11426_/Q _09154_/X _09163_/X vssd1 vssd1 vccd1 vccd1 _11426_/D sky130_fd_sc_hd__a21o_1
XFILLER_33_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06376_ _11322_/Q _06738_/A2 _06739_/A2 _11294_/Q vssd1 vssd1 vccd1 vccd1 _06376_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08115_ _10884_/Q _10132_/A0 _08120_/S vssd1 vssd1 vccd1 vccd1 _08116_/B sky130_fd_sc_hd__mux2_1
X_05327_ _10458_/Q _10457_/Q _06967_/A vssd1 vssd1 vccd1 vccd1 _05329_/C sky130_fd_sc_hd__mux2_1
XFILLER_147_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09095_ _11395_/Q _09099_/B vssd1 vssd1 vccd1 vccd1 _09095_/X sky130_fd_sc_hd__or2_1
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_2__f_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_2__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_08046_ _10849_/Q _10132_/A0 _08051_/S vssd1 vssd1 vccd1 vccd1 _08047_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05258_ _05258_/A _05258_/B _05258_/C _05258_/D vssd1 vssd1 vccd1 vccd1 _05259_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05189_ _05189_/A _05189_/B _05189_/C _05189_/D vssd1 vssd1 vccd1 vccd1 _05190_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_153_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09997_ _11685_/Q _09977_/X _09996_/X vssd1 vssd1 vccd1 vccd1 _11685_/D sky130_fd_sc_hd__a21o_1
XFILLER_153_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08948_ _09538_/A _09538_/B vssd1 vssd1 vccd1 vccd1 _09668_/D sky130_fd_sc_hd__nand2_2
XFILLER_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ _08931_/A1 _08890_/S _08878_/X _09078_/C1 vssd1 vssd1 vccd1 vccd1 _11296_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ _11777_/CLK _10910_/D vssd1 vssd1 vccd1 vccd1 _10910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ _11280_/CLK _10841_/D vssd1 vssd1 vccd1 vccd1 _10841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ _11471_/CLK _10772_/D vssd1 vssd1 vccd1 vccd1 _10772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11324_ _11385_/CLK _11324_/D vssd1 vssd1 vccd1 vccd1 _11324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11255_ _11572_/CLK _11255_/D vssd1 vssd1 vccd1 vccd1 _11255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10206_ _11809_/CLK _10206_/D vssd1 vssd1 vccd1 vccd1 _10206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11186_ _11186_/CLK _11186_/D vssd1 vssd1 vccd1 vccd1 _11186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10137_ _10137_/A _10137_/B _10159_/C vssd1 vssd1 vccd1 vccd1 _10137_/X sky130_fd_sc_hd__or3_4
XFILLER_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ _10115_/A0 _11729_/Q _10071_/S vssd1 vssd1 vccd1 vccd1 _11729_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06230_ _10263_/Q _06230_/A2 _06540_/B1 _10200_/Q vssd1 vssd1 vccd1 vccd1 _06230_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06161_ _10648_/Q _06161_/A2 _06159_/X _06160_/X vssd1 vssd1 vccd1 vccd1 _06161_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05112_ _05112_/A _05112_/B _05112_/C _05112_/D vssd1 vssd1 vccd1 vccd1 _05113_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06092_ _11384_/Q _09060_/A _06088_/X _06091_/X vssd1 vssd1 vccd1 vccd1 _06093_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_89_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09920_ _10488_/Q _09570_/B _09572_/C _10494_/Q _09919_/X vssd1 vssd1 vccd1 vccd1
+ _09925_/B sky130_fd_sc_hd__a221o_1
XFILLER_116_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout706 _10087_/C vssd1 vssd1 vccd1 vccd1 _10159_/C sky130_fd_sc_hd__clkbuf_8
Xfanout717 _06105_/B1 vssd1 vssd1 vccd1 vccd1 _07819_/A sky130_fd_sc_hd__clkbuf_16
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09851_ _09908_/A _09851_/B vssd1 vssd1 vccd1 vccd1 _09851_/Y sky130_fd_sc_hd__nor2_2
Xfanout728 fanout738/X vssd1 vssd1 vccd1 vccd1 _06871_/B1 sky130_fd_sc_hd__buf_4
XFILLER_59_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _09292_/A vssd1 vssd1 vccd1 vccd1 _08286_/A sky130_fd_sc_hd__buf_12
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08802_ _08893_/A1 _11257_/Q _08802_/S vssd1 vssd1 vccd1 vccd1 _08803_/B sky130_fd_sc_hd__mux2_1
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _11648_/Q _08950_/B _09781_/X _09407_/A vssd1 vssd1 vccd1 vccd1 _11648_/D
+ sky130_fd_sc_hd__o211a_1
X_06994_ _10264_/Q _06976_/X _06993_/X vssd1 vssd1 vccd1 vccd1 _10264_/D sky130_fd_sc_hd__a21o_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _08733_/A _08733_/B vssd1 vssd1 vccd1 vccd1 _11223_/D sky130_fd_sc_hd__or2_1
XFILLER_22_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05945_ _05095_/Y _05907_/X _05918_/X _05923_/X vssd1 vssd1 vccd1 vccd1 _05945_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08664_ _08664_/A _08664_/B vssd1 vssd1 vccd1 vccd1 _11187_/D sky130_fd_sc_hd__or2_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05876_ _10870_/Q _06415_/A2 _06453_/B1 _10986_/Q vssd1 vssd1 vccd1 vccd1 _05876_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ _10591_/Q _07613_/Y _07614_/Y _07324_/X vssd1 vssd1 vccd1 vccd1 _10591_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _09111_/A1 _11152_/Q _08623_/S vssd1 vssd1 vccd1 vccd1 _08596_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07546_ _08536_/A _07546_/B vssd1 vssd1 vccd1 vccd1 _10556_/D sky130_fd_sc_hd__or2_1
XFILLER_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07477_ _10047_/A1 _10517_/Q _07477_/S vssd1 vssd1 vccd1 vccd1 _07478_/B sky130_fd_sc_hd__mux2_1
X_09216_ _09216_/A0 _11457_/Q _09218_/S vssd1 vssd1 vccd1 vccd1 _09216_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06428_ _10883_/Q _06468_/B _06641_/A2 _10614_/Q _06427_/X vssd1 vssd1 vccd1 vccd1
+ _06428_/X sky130_fd_sc_hd__o221a_1
XFILLER_155_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09147_ _10175_/A1 _09149_/B _10166_/B1 vssd1 vssd1 vccd1 vccd1 _09147_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06359_ _11527_/Q _09326_/A _09977_/A _11685_/Q vssd1 vssd1 vccd1 vccd1 _06359_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09078_ _09172_/A1 _09060_/X _09077_/X _09078_/C1 vssd1 vssd1 vccd1 vccd1 _11387_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ _10839_/Q _08037_/B vssd1 vssd1 vccd1 vccd1 _08029_/X sky130_fd_sc_hd__or2_1
XFILLER_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11040_ _11329_/CLK _11040_/D vssd1 vssd1 vccd1 vccd1 _11040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11873_ input86/X vssd1 vssd1 vccd1 vccd1 _11873_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _11270_/CLK _10824_/D vssd1 vssd1 vccd1 vccd1 _10824_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10755_ _11573_/CLK _10755_/D vssd1 vssd1 vccd1 vccd1 _10755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10686_ _11703_/CLK _10686_/D vssd1 vssd1 vccd1 vccd1 _10686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _11307_/CLK _11307_/D vssd1 vssd1 vccd1 vccd1 _11307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11238_ _11485_/CLK _11238_/D vssd1 vssd1 vccd1 vccd1 _11238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11169_ _11812_/CLK _11169_/D vssd1 vssd1 vccd1 vccd1 _11169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05730_ input78/X _10255_/D vssd1 vssd1 vccd1 vccd1 _05730_/Y sky130_fd_sc_hd__nand2_8
XFILLER_110_1347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05661_ _05661_/A _05661_/B _05661_/C _05661_/D vssd1 vssd1 vccd1 vccd1 _05668_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07400_ _10026_/A _07400_/B vssd1 vssd1 vccd1 vccd1 _10476_/D sky130_fd_sc_hd__or2_1
XFILLER_17_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08380_ _08380_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08380_/Y sky130_fd_sc_hd__nand2_1
X_05592_ _05628_/A2 _11485_/Q _11482_/Q _05628_/B1 vssd1 vssd1 vccd1 vccd1 _05592_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07331_ _10431_/Q _07322_/Y _07326_/Y _07316_/X vssd1 vssd1 vccd1 vccd1 _10431_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07262_ _07936_/A _07262_/B vssd1 vssd1 vccd1 vccd1 _10399_/D sky130_fd_sc_hd__or2_1
XFILLER_143_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09001_ _09256_/A1 _09013_/B _08761_/A vssd1 vssd1 vccd1 vccd1 _09001_/X sky130_fd_sc_hd__a21o_1
X_06213_ _11525_/Q _08383_/A _08245_/A _11485_/Q vssd1 vssd1 vccd1 vccd1 _06213_/X
+ sky130_fd_sc_hd__o22a_1
X_07193_ _07333_/B _07191_/B _07192_/A _10356_/Q _07333_/A vssd1 vssd1 vccd1 vccd1
+ _10356_/D sky130_fd_sc_hd__a221o_1
XFILLER_118_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06144_ _07082_/A _06142_/X _06143_/X _05816_/A vssd1 vssd1 vccd1 vccd1 _06144_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_118_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06075_ _06633_/A _06075_/B _06075_/C vssd1 vssd1 vccd1 vccd1 _06075_/X sky130_fd_sc_hd__or3_1
XFILLER_133_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09903_ _11708_/Q _09568_/C _09944_/B1 _11710_/Q vssd1 vssd1 vccd1 vccd1 _09903_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout503 _09122_/C1 vssd1 vssd1 vccd1 vccd1 _09078_/C1 sky130_fd_sc_hd__buf_4
XFILLER_154_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout514 _08050_/A vssd1 vssd1 vccd1 vccd1 _08196_/A sky130_fd_sc_hd__buf_4
Xfanout525 fanout536/X vssd1 vssd1 vccd1 vccd1 _07659_/A sky130_fd_sc_hd__buf_4
XFILLER_98_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout536 _06898_/Y vssd1 vssd1 vccd1 vccd1 fanout536/X sky130_fd_sc_hd__buf_6
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout547 _07812_/A vssd1 vssd1 vccd1 vccd1 _07922_/A sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_127_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10798_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09834_ _11453_/Q _09886_/A2 _09876_/B1 _10774_/Q vssd1 vssd1 vccd1 vccd1 _09834_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout558 _08618_/A vssd1 vssd1 vccd1 vccd1 _08851_/A sky130_fd_sc_hd__buf_4
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout569 _08670_/A vssd1 vssd1 vccd1 vccd1 _08941_/A sky130_fd_sc_hd__clkbuf_4
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09765_ _09522_/B _09722_/Y _09758_/Y _06962_/X vssd1 vssd1 vccd1 vccd1 _09765_/X
+ sky130_fd_sc_hd__a22o_1
X_06977_ _10256_/Q _06995_/B vssd1 vssd1 vccd1 vccd1 _06977_/X sky130_fd_sc_hd__or2_1
XFILLER_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08716_ _08810_/A _08716_/B vssd1 vssd1 vccd1 vccd1 _11213_/D sky130_fd_sc_hd__or2_1
XFILLER_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05928_ _11305_/Q _10010_/A _05924_/X _05927_/X vssd1 vssd1 vccd1 vccd1 _05934_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09696_ _11635_/Q _11639_/Q _09702_/S vssd1 vssd1 vccd1 vccd1 _09697_/B sky130_fd_sc_hd__mux2_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08647_ _08647_/A _08647_/B _10119_/B _10119_/C vssd1 vssd1 vccd1 vccd1 _08647_/X
+ sky130_fd_sc_hd__or4_2
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05859_ _11104_/Q _06716_/A2 _05855_/X _05858_/X vssd1 vssd1 vccd1 vccd1 _05859_/X
+ sky130_fd_sc_hd__o211a_4
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ _08578_/A _08578_/B vssd1 vssd1 vccd1 vccd1 _11144_/D sky130_fd_sc_hd__and2_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ _10051_/A1 _10549_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _07530_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10540_ _11472_/CLK _10540_/D vssd1 vssd1 vccd1 vccd1 _10540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10471_ _11136_/CLK _10471_/D vssd1 vssd1 vccd1 vccd1 _10471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11023_ _11023_/CLK _11023_/D vssd1 vssd1 vccd1 vccd1 _11023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ _11462_/CLK _10807_/D vssd1 vssd1 vccd1 vccd1 _10807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11787_ _11791_/CLK _11787_/D vssd1 vssd1 vccd1 vccd1 _11787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10738_ _11768_/CLK _10738_/D vssd1 vssd1 vccd1 vccd1 _10738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10669_ _10773_/CLK _10669_/D vssd1 vssd1 vccd1 vccd1 _10669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput128 _11812_/Q vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_4
Xoutput139 _11619_/Q vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__buf_4
XFILLER_126_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06900_ _06900_/A _07151_/C _07151_/D vssd1 vssd1 vccd1 vccd1 _09270_/B sky130_fd_sc_hd__and3_4
XFILLER_110_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07880_ _07025_/A _07890_/A2 _07879_/X _07932_/C1 vssd1 vssd1 vccd1 vccd1 _10758_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06831_ _10395_/Q _06860_/A2 _06827_/X _06830_/X vssd1 vssd1 vccd1 vccd1 _06831_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09550_ _05076_/A _09541_/Y _09549_/X _09833_/A vssd1 vssd1 vccd1 vccd1 _11627_/D
+ sky130_fd_sc_hd__o211a_1
X_06762_ _10548_/Q _07440_/A vssd1 vssd1 vccd1 vccd1 _06762_/X sky130_fd_sc_hd__or2_1
XFILLER_23_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08501_ _08760_/A0 _11101_/Q _08501_/S vssd1 vssd1 vccd1 vccd1 _08502_/B sky130_fd_sc_hd__mux2_1
XFILLER_110_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05713_ _11049_/Q _05579_/Y _05597_/Y _11040_/Q vssd1 vssd1 vccd1 vccd1 _05713_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09481_ _11604_/Q _09554_/A vssd1 vssd1 vccd1 vccd1 _09481_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06693_ _10670_/Q _06875_/B1 _06692_/X _06808_/C1 vssd1 vssd1 vccd1 vccd1 _06693_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08432_ _11057_/Q _08425_/Y _08426_/Y _07093_/X vssd1 vssd1 vccd1 vccd1 _11057_/D
+ sky130_fd_sc_hd__o22a_1
X_05644_ _05644_/A _05644_/B _05644_/C vssd1 vssd1 vccd1 vccd1 _05644_/X sky130_fd_sc_hd__or3_4
X_08363_ _08469_/A _08360_/S _08362_/X _09022_/C1 vssd1 vssd1 vccd1 vccd1 _11024_/D
+ sky130_fd_sc_hd__o211a_1
X_05575_ _05629_/A2 _11367_/Q _11361_/Q _05629_/B1 vssd1 vssd1 vccd1 vccd1 _05575_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07314_ _08902_/B _07314_/B vssd1 vssd1 vccd1 vccd1 _07314_/X sky130_fd_sc_hd__or2_4
X_08294_ _10980_/Q _07617_/X _08298_/S vssd1 vssd1 vccd1 vccd1 _10980_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07245_ _07309_/A _07245_/B vssd1 vssd1 vccd1 vccd1 _07245_/X sky130_fd_sc_hd__or2_1
XFILLER_30_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07176_ _10349_/Q _09228_/B vssd1 vssd1 vccd1 vccd1 _07176_/X sky130_fd_sc_hd__or2_1
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06127_ _11128_/Q _06635_/A2 _08647_/B _11177_/Q _06126_/X vssd1 vssd1 vccd1 vccd1
+ _06127_/X sky130_fd_sc_hd__o221a_1
XFILLER_106_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06058_ _11259_/Q _06514_/A2 _05865_/B _11770_/Q _06057_/X vssd1 vssd1 vccd1 vccd1
+ _06059_/B sky130_fd_sc_hd__o221a_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout300 _07623_/X vssd1 vssd1 vccd1 vccd1 _08459_/S sky130_fd_sc_hd__buf_4
Xfanout311 _07752_/B vssd1 vssd1 vccd1 vccd1 _07754_/B sky130_fd_sc_hd__buf_6
XFILLER_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout322 _07259_/S vssd1 vssd1 vccd1 vccd1 _07277_/S sky130_fd_sc_hd__clkbuf_4
Xfanout333 _07150_/A2 vssd1 vssd1 vccd1 vccd1 _07135_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout344 _07225_/X vssd1 vssd1 vccd1 vccd1 _08441_/B2 sky130_fd_sc_hd__buf_12
XFILLER_86_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout355 _10010_/B vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__buf_12
XFILLER_101_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout366 _07052_/X vssd1 vssd1 vccd1 vccd1 _07617_/B sky130_fd_sc_hd__buf_8
XFILLER_101_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09817_ _11643_/Q _09817_/B vssd1 vssd1 vccd1 vccd1 _09817_/Y sky130_fd_sc_hd__xnor2_2
Xfanout377 _08322_/A vssd1 vssd1 vccd1 vccd1 _08902_/B sky130_fd_sc_hd__buf_12
Xfanout388 _07004_/Y vssd1 vssd1 vccd1 vccd1 _07614_/A sky130_fd_sc_hd__buf_6
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout399 _05434_/Y vssd1 vssd1 vccd1 vccd1 _09877_/B1 sky130_fd_sc_hd__buf_4
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09748_ _10540_/Q _09573_/A _09872_/A2 _10550_/Q _09747_/X vssd1 vssd1 vccd1 vccd1
+ _09749_/D sky130_fd_sc_hd__a221o_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _11602_/Q _09679_/B vssd1 vssd1 vccd1 vccd1 _09681_/C sky130_fd_sc_hd__nand2_1
XFILLER_76_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11710_/CLK _11710_/D vssd1 vssd1 vccd1 vccd1 _11710_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_95_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _10804_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11269_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11641_ _11641_/CLK _11641_/D vssd1 vssd1 vccd1 vccd1 _11641_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11572_ _11572_/CLK _11572_/D vssd1 vssd1 vccd1 vccd1 _11572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10523_ _11308_/CLK _10523_/D vssd1 vssd1 vccd1 vccd1 _10523_/Q sky130_fd_sc_hd__dfxtp_2
Xinput19 rom_value[18] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10454_ _11776_/CLK _10454_/D vssd1 vssd1 vccd1 vccd1 _10454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10385_ _11133_/CLK _10385_/D vssd1 vssd1 vccd1 vccd1 _10385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11006_ _11235_/CLK _11006_/D vssd1 vssd1 vccd1 vccd1 _11006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05360_ _10988_/Q _10987_/Q _05429_/S vssd1 vssd1 vccd1 vccd1 _05362_/C sky130_fd_sc_hd__mux2_1
XFILLER_144_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05291_ _05291_/A _05291_/B _05291_/C _05291_/D vssd1 vssd1 vccd1 vccd1 _05291_/Y
+ sky130_fd_sc_hd__nor4_4
X_07030_ _10274_/Q _07029_/X _07044_/S vssd1 vssd1 vccd1 vccd1 _10274_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08981_ _11343_/Q _08989_/B vssd1 vssd1 vccd1 vccd1 _08981_/X sky130_fd_sc_hd__or2_1
XFILLER_64_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07932_ _07932_/A1 _09218_/S _07931_/X _07932_/C1 vssd1 vssd1 vccd1 vccd1 _10783_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07863_ _10750_/Q _07883_/B vssd1 vssd1 vccd1 vccd1 _07863_/X sky130_fd_sc_hd__or2_1
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09602_ _10385_/Q _09568_/C _09948_/B1 _10386_/Q vssd1 vssd1 vccd1 vccd1 _09617_/A
+ sky130_fd_sc_hd__a22o_2
X_06814_ _11446_/Q _07777_/A _07254_/A _11439_/Q vssd1 vssd1 vccd1 vccd1 _06814_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_83_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07794_ _07796_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _10704_/D sky130_fd_sc_hd__or2_1
X_09533_ _09528_/A _09502_/B _09508_/Y _09532_/X _09529_/A vssd1 vssd1 vccd1 vccd1
+ _11621_/D sky130_fd_sc_hd__o311a_1
X_06745_ _10627_/Q _06860_/A2 _06710_/B _10731_/Q vssd1 vssd1 vccd1 vccd1 _06745_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09464_ input37/X input14/X input23/X input31/X _11576_/Q _11577_/Q vssd1 vssd1 vccd1
+ vccd1 _09464_/X sky130_fd_sc_hd__mux4_1
X_06676_ _06670_/X _06675_/X _06743_/B vssd1 vssd1 vccd1 vccd1 _06676_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08415_ _08684_/A _08415_/B vssd1 vssd1 vccd1 vccd1 _11048_/D sky130_fd_sc_hd__or2_1
X_05627_ _05627_/A _05627_/B vssd1 vssd1 vccd1 vccd1 _05627_/Y sky130_fd_sc_hd__nor2_8
X_09395_ _09395_/A0 _11561_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _11561_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08346_ _10114_/A0 _11016_/Q _08354_/S vssd1 vssd1 vccd1 vccd1 _08347_/B sky130_fd_sc_hd__mux2_1
X_05558_ _05618_/A1 _11342_/Q _11339_/Q _05606_/B2 _05556_/X vssd1 vssd1 vccd1 vccd1
+ _05561_/A sky130_fd_sc_hd__a221o_4
XFILLER_123_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08277_ _08684_/A _08277_/B vssd1 vssd1 vccd1 vccd1 _10970_/D sky130_fd_sc_hd__or2_1
X_05489_ _10234_/Q input45/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05489_/X sky130_fd_sc_hd__mux2_1
X_07228_ _07227_/X _10381_/Q _07249_/S vssd1 vssd1 vccd1 vccd1 _10381_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_142_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11781_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07159_ _07790_/A _07159_/B vssd1 vssd1 vccd1 vccd1 _10340_/D sky130_fd_sc_hd__or2_1
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10170_ _11797_/Q _10176_/B vssd1 vssd1 vccd1 vccd1 _10170_/X sky130_fd_sc_hd__or2_1
XFILLER_121_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _11812_/CLK _11624_/D vssd1 vssd1 vccd1 vccd1 _11624_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_156_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11555_ _11763_/CLK _11555_/D vssd1 vssd1 vccd1 vccd1 _11555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10506_ _11462_/CLK _10506_/D vssd1 vssd1 vccd1 vccd1 _10506_/Q sky130_fd_sc_hd__dfxtp_1
X_11486_ _11809_/CLK _11486_/D vssd1 vssd1 vccd1 vccd1 _11486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10437_ _11768_/CLK _10437_/D vssd1 vssd1 vccd1 vccd1 _10437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10368_ _10727_/CLK _10368_/D vssd1 vssd1 vccd1 vccd1 _10368_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _11745_/CLK _10299_/D vssd1 vssd1 vccd1 vccd1 _10299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06530_ _11201_/Q _06645_/A2 _09109_/A _11251_/Q vssd1 vssd1 vccd1 vccd1 _06530_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06461_ _10896_/Q _08123_/A _06457_/X _06460_/X vssd1 vssd1 vccd1 vccd1 _06461_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_34_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08200_ _08200_/A _10119_/B _09038_/C vssd1 vssd1 vccd1 vccd1 _08200_/X sky130_fd_sc_hd__or3_2
XFILLER_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05412_ _05412_/A _05412_/B vssd1 vssd1 vccd1 vccd1 _05412_/Y sky130_fd_sc_hd__nor2_4
X_09180_ _11434_/Q _07613_/A _09175_/B _09179_/X vssd1 vssd1 vccd1 vccd1 _11434_/D
+ sky130_fd_sc_hd__o31a_1
X_06392_ _11018_/Q _06630_/B1 _06391_/X _06392_/C1 vssd1 vssd1 vccd1 vccd1 _06392_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08131_ _09396_/A0 _08140_/S _08130_/X _08345_/C1 vssd1 vssd1 vccd1 vccd1 _10891_/D
+ sky130_fd_sc_hd__o211a_1
X_05343_ _11102_/Q _11101_/Q _05471_/A vssd1 vssd1 vccd1 vccd1 _05345_/C sky130_fd_sc_hd__mux2_1
XFILLER_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08062_ _08590_/A _08062_/B vssd1 vssd1 vccd1 vccd1 _10856_/D sky130_fd_sc_hd__or2_1
X_05274_ _10813_/Q _10812_/Q _05372_/S vssd1 vssd1 vccd1 vccd1 _05275_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_4_1__f_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_146_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07013_ _07227_/B _07318_/A vssd1 vssd1 vccd1 vccd1 _07013_/X sky130_fd_sc_hd__or2_4
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08964_ _08963_/X _11334_/Q _09830_/B vssd1 vssd1 vccd1 vccd1 _08965_/B sky130_fd_sc_hd__mux2_1
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07915_ _08931_/A1 _10775_/Q _09218_/S vssd1 vssd1 vccd1 vccd1 _07916_/B sky130_fd_sc_hd__mux2_1
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08895_ _08947_/A1 _08874_/S _08894_/X _08947_/C1 vssd1 vssd1 vccd1 vccd1 _11304_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07846_ _07235_/X _10741_/Q _07846_/S vssd1 vssd1 vccd1 vccd1 _10741_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07777_ _07777_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _09192_/B sky130_fd_sc_hd__nor2_2
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06728_ _10573_/Q _06877_/B1 _06728_/B1 _10546_/Q vssd1 vssd1 vccd1 vccd1 _06728_/X
+ sky130_fd_sc_hd__o22a_1
X_09516_ _09516_/A vssd1 vssd1 vccd1 vccd1 _09516_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09447_ _09539_/A _09447_/B vssd1 vssd1 vccd1 vccd1 _09447_/Y sky130_fd_sc_hd__nand2_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06659_ _11118_/Q _09081_/A _06657_/X _06658_/X vssd1 vssd1 vccd1 vccd1 _06659_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ _10106_/A1 _09376_/B _10156_/B1 vssd1 vssd1 vccd1 vccd1 _09378_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ _11004_/Q _08322_/Y _08325_/Y _07019_/X vssd1 vssd1 vccd1 vccd1 _11004_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11340_ _11495_/CLK _11340_/D vssd1 vssd1 vccd1 vccd1 _11340_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11271_ _11601_/CLK _11271_/D vssd1 vssd1 vccd1 vccd1 _11271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10222_ _11307_/CLK _10222_/D vssd1 vssd1 vccd1 vccd1 _10222_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _10153_/A1 _10137_/X _10152_/X _10153_/C1 vssd1 vssd1 vccd1 vccd1 _11789_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10084_ _11744_/Q _07451_/X _10085_/S vssd1 vssd1 vccd1 vccd1 _11744_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10986_ _11633_/CLK _10986_/D vssd1 vssd1 vccd1 vccd1 _10986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ _11607_/CLK _11607_/D vssd1 vssd1 vccd1 vccd1 _11607_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11538_ _11801_/CLK _11538_/D vssd1 vssd1 vccd1 vccd1 _11538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11469_ _11471_/CLK _11469_/D vssd1 vssd1 vccd1 vccd1 _11469_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05961_ _11372_/Q _06221_/A2 _05957_/X _05960_/X vssd1 vssd1 vccd1 vccd1 _05962_/C
+ sky130_fd_sc_hd__o211a_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07700_ _10648_/Q _07693_/Y _07697_/Y _07016_/X vssd1 vssd1 vccd1 vccd1 _10648_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08680_ _08941_/A _08680_/B vssd1 vssd1 vccd1 vccd1 _11194_/D sky130_fd_sc_hd__or2_1
X_05892_ _11424_/Q _08668_/A _09038_/A _11371_/Q vssd1 vssd1 vccd1 vccd1 _05892_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07631_ _08816_/A _08820_/S vssd1 vssd1 vccd1 vccd1 _07637_/S sky130_fd_sc_hd__or2_4
XFILLER_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07562_ _08781_/A _07562_/B vssd1 vssd1 vccd1 vccd1 _10564_/D sky130_fd_sc_hd__or2_1
XFILLER_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ _11501_/Q _09293_/X _09300_/X vssd1 vssd1 vccd1 vccd1 _11501_/D sky130_fd_sc_hd__a21o_1
X_06513_ _10445_/Q _06513_/A2 _06636_/A2 _11079_/Q _06550_/C1 vssd1 vssd1 vccd1 vccd1
+ _06513_/X sky130_fd_sc_hd__o221a_1
XFILLER_80_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07493_ _10529_/Q _07496_/S _07141_/X _07078_/B _07451_/A vssd1 vssd1 vccd1 vccd1
+ _10529_/D sky130_fd_sc_hd__a221o_1
XFILLER_107_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09232_ _11466_/Q _09226_/Y _09229_/Y _09232_/B2 vssd1 vssd1 vccd1 vccd1 _11466_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06444_ _11323_/Q _06648_/A2 _09131_/A _11295_/Q _08243_/B vssd1 vssd1 vccd1 vccd1
+ _06444_/X sky130_fd_sc_hd__a221o_1
XFILLER_142_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09163_ _10168_/A1 _09171_/B _10166_/B1 vssd1 vssd1 vccd1 vccd1 _09163_/X sky130_fd_sc_hd__a21o_1
X_06375_ _06365_/X _06366_/X _06369_/X _06374_/X vssd1 vssd1 vccd1 vccd1 _06375_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08114_ _10883_/Q _08102_/S _07642_/S _07316_/B vssd1 vssd1 vccd1 vccd1 _10883_/D
+ sky130_fd_sc_hd__o22a_1
X_05326_ _10845_/Q _10844_/Q _05326_/S vssd1 vssd1 vccd1 vccd1 _05329_/B sky130_fd_sc_hd__mux2_1
X_09094_ _11394_/Q _09082_/X _09093_/X vssd1 vssd1 vccd1 vccd1 _11394_/D sky130_fd_sc_hd__a21o_1
XFILLER_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08045_ _10848_/Q _07364_/X _07365_/Y _07316_/B vssd1 vssd1 vccd1 vccd1 _10848_/D
+ sky130_fd_sc_hd__o22a_1
X_05257_ _11086_/Q _11085_/Q _05399_/S vssd1 vssd1 vccd1 vccd1 _05258_/D sky130_fd_sc_hd__mux2_2
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05188_ _10839_/Q _10838_/Q _06945_/B vssd1 vssd1 vccd1 vccd1 _05189_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09996_ _10178_/A1 _09994_/B _08851_/A vssd1 vssd1 vccd1 vccd1 _09996_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08947_ _08947_/A1 _08907_/X _08946_/X _08947_/C1 vssd1 vssd1 vccd1 vccd1 _11332_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08878_ _11296_/Q _08894_/B vssd1 vssd1 vccd1 vccd1 _08878_/X sky130_fd_sc_hd__or2_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07829_ _07061_/A _07820_/B _07956_/S _10724_/Q vssd1 vssd1 vccd1 vccd1 _10724_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10840_ _11657_/CLK _10840_/D vssd1 vssd1 vccd1 vccd1 _10840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10771_ _11644_/CLK _10771_/D vssd1 vssd1 vccd1 vccd1 _10771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11323_ _11332_/CLK _11323_/D vssd1 vssd1 vccd1 vccd1 _11323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11254_ _11329_/CLK _11254_/D vssd1 vssd1 vccd1 vccd1 _11254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _11810_/CLK _10205_/D vssd1 vssd1 vccd1 vccd1 _10205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11185_ _11186_/CLK _11185_/D vssd1 vssd1 vccd1 vccd1 _11185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10136_ _10136_/A _10136_/B _10136_/C vssd1 vssd1 vccd1 vccd1 _10154_/B sky130_fd_sc_hd__and3_4
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10067_ _10114_/A0 _11728_/Q _10071_/S vssd1 vssd1 vccd1 vccd1 _11728_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10969_ _11575_/CLK _10969_/D vssd1 vssd1 vccd1 vccd1 _10969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06160_ _11311_/Q _06459_/A2 _06459_/B1 _10873_/Q vssd1 vssd1 vccd1 vccd1 _06160_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05111_ _11268_/Q _11267_/Q _09430_/B vssd1 vssd1 vccd1 vccd1 _05112_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06091_ _11427_/Q _08668_/A _06090_/X _06670_/D1 vssd1 vssd1 vccd1 vccd1 _06091_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ _09850_/A _09850_/B _09850_/C _09850_/D vssd1 vssd1 vccd1 vccd1 _09851_/B
+ sky130_fd_sc_hd__or4_4
Xfanout707 _07298_/X vssd1 vssd1 vccd1 vccd1 _10087_/C sky130_fd_sc_hd__buf_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout718 _06105_/B1 vssd1 vssd1 vccd1 vccd1 _07827_/A2 sky130_fd_sc_hd__buf_4
Xfanout729 _06728_/B1 vssd1 vssd1 vccd1 vccd1 _07440_/A sky130_fd_sc_hd__buf_8
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08801_ _09237_/A0 _08792_/S _08800_/X _07003_/B vssd1 vssd1 vccd1 vccd1 _11256_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06993_ _10105_/A1 _06995_/B _08664_/A vssd1 vssd1 vccd1 vccd1 _06993_/X sky130_fd_sc_hd__a21o_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _11647_/Q _09404_/Y _09780_/X _09681_/B vssd1 vssd1 vccd1 vccd1 _09781_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _07092_/A _11223_/Q _08742_/S vssd1 vssd1 vccd1 vccd1 _08733_/B sky130_fd_sc_hd__mux2_1
X_05944_ _11089_/Q _06589_/A2 _05940_/X _05943_/X vssd1 vssd1 vccd1 vccd1 _05944_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08663_ _11187_/Q _08760_/A0 _08663_/S vssd1 vssd1 vccd1 vccd1 _08664_/B sky130_fd_sc_hd__mux2_1
X_05875_ _11062_/Q _06629_/A2 _05871_/X _05874_/X vssd1 vssd1 vccd1 vccd1 _05875_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07614_ _07614_/A _08035_/S vssd1 vssd1 vccd1 vccd1 _07614_/Y sky130_fd_sc_hd__nand2_2
XFILLER_42_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08594_ _08594_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08594_/X sky130_fd_sc_hd__or2_4
XFILLER_35_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07545_ _10015_/A0 _10556_/Q _07591_/S vssd1 vssd1 vccd1 vccd1 _07546_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07476_ _07476_/A _07476_/B vssd1 vssd1 vccd1 vccd1 _10516_/D sky130_fd_sc_hd__or2_1
XFILLER_22_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06427_ _11227_/Q _08650_/A _06639_/B1 _10453_/Q vssd1 vssd1 vccd1 vccd1 _06427_/X
+ sky130_fd_sc_hd__o22a_1
X_09215_ _11456_/Q _09206_/Y _09214_/X _09229_/A vssd1 vssd1 vccd1 vccd1 _11456_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09146_ _10172_/A1 _09132_/X _09145_/X _10175_/C1 vssd1 vssd1 vccd1 vccd1 _11418_/D
+ sky130_fd_sc_hd__o211a_1
X_06358_ _11421_/Q _06718_/B1 _06354_/X _06357_/X vssd1 vssd1 vccd1 vccd1 _06364_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_147_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05309_ _11022_/Q _11021_/Q _09680_/C vssd1 vssd1 vccd1 vccd1 _05312_/B sky130_fd_sc_hd__mux2_1
X_09077_ _11387_/Q _09077_/B vssd1 vssd1 vccd1 vccd1 _09077_/X sky130_fd_sc_hd__or2_1
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06289_ _08243_/A _11872_/A vssd1 vssd1 vccd1 vccd1 _06901_/A sky130_fd_sc_hd__nand2_1
XFILLER_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_49_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11366_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08028_ _08847_/A _08028_/B vssd1 vssd1 vccd1 vccd1 _10838_/D sky130_fd_sc_hd__or2_1
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09979_ _11676_/Q _09977_/X _09978_/X vssd1 vssd1 vccd1 vccd1 _11676_/D sky130_fd_sc_hd__a21o_1
XFILLER_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11872_/A vssd1 vssd1 vccd1 vccd1 _11872_/X sky130_fd_sc_hd__buf_2
XFILLER_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ _11634_/CLK _10823_/D vssd1 vssd1 vccd1 vccd1 _10823_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ _11622_/CLK _10754_/D vssd1 vssd1 vccd1 vccd1 _10754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10685_ _10798_/CLK _10685_/D vssd1 vssd1 vccd1 vccd1 _10685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11306_ _11776_/CLK _11306_/D vssd1 vssd1 vccd1 vccd1 _11306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11237_ _11366_/CLK _11237_/D vssd1 vssd1 vccd1 vccd1 _11237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11168_ _11572_/CLK _11168_/D vssd1 vssd1 vccd1 vccd1 _11168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10119_ _10119_/A _10119_/B _10119_/C vssd1 vssd1 vccd1 vccd1 _10119_/X sky130_fd_sc_hd__or3_2
X_11099_ _11151_/CLK _11099_/D vssd1 vssd1 vccd1 vccd1 _11099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05660_ _11241_/Q _05531_/Y _05555_/Y _11250_/Q vssd1 vssd1 vccd1 vccd1 _05661_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05591_ _05591_/A _05591_/B vssd1 vssd1 vccd1 vccd1 _05591_/Y sky130_fd_sc_hd__nor2_8
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07330_ _10430_/Q _07322_/Y _07326_/Y _07019_/X vssd1 vssd1 vccd1 vccd1 _10430_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07261_ _10019_/A0 _10399_/Q _09184_/S vssd1 vssd1 vccd1 vccd1 _07262_/B sky130_fd_sc_hd__mux2_1
XFILLER_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09000_ _10183_/A0 _08994_/X _08999_/X _09036_/C1 vssd1 vssd1 vccd1 vccd1 _11351_/D
+ sky130_fd_sc_hd__o211a_1
X_06212_ _06450_/A _10229_/Q vssd1 vssd1 vccd1 vccd1 _06212_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07192_ _07192_/A vssd1 vssd1 vccd1 vccd1 _07192_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06143_ _06633_/A _06136_/X _06141_/X _07081_/A _06131_/X vssd1 vssd1 vccd1 vccd1
+ _06143_/X sky130_fd_sc_hd__o311a_2
XFILLER_133_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06074_ _11091_/Q _06629_/B1 _06070_/X _06073_/X vssd1 vssd1 vccd1 vccd1 _06075_/C
+ sky130_fd_sc_hd__o211a_1
X_09902_ _11697_/Q _09568_/D _09571_/D _11700_/Q _09901_/X vssd1 vssd1 vccd1 vccd1
+ _09907_/B sky130_fd_sc_hd__a221o_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout504 _09122_/C1 vssd1 vssd1 vccd1 vccd1 _09289_/C1 sky130_fd_sc_hd__buf_4
Xfanout515 _08050_/A vssd1 vssd1 vccd1 vccd1 _08749_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout526 _08835_/A vssd1 vssd1 vccd1 vccd1 _08839_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout537 _10056_/A vssd1 vssd1 vccd1 vccd1 _10058_/A sky130_fd_sc_hd__clkbuf_4
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _09833_/A _09833_/B vssd1 vssd1 vccd1 vccd1 _11657_/D sky130_fd_sc_hd__and2_1
XFILLER_98_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout548 fanout555/X vssd1 vssd1 vccd1 vccd1 _07812_/A sky130_fd_sc_hd__buf_2
XFILLER_150_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout559 _08618_/A vssd1 vssd1 vccd1 vccd1 _10178_/B1 sky130_fd_sc_hd__clkbuf_8
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _11644_/Q _09763_/X _09770_/S vssd1 vssd1 vccd1 vccd1 _11644_/D sky130_fd_sc_hd__mux2_1
X_06976_ _06976_/A _10180_/C _10137_/B vssd1 vssd1 vccd1 vccd1 _06976_/X sky130_fd_sc_hd__or3_4
XFILLER_100_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08715_ _11213_/Q _07015_/A _08726_/S vssd1 vssd1 vccd1 vccd1 _08716_/B sky130_fd_sc_hd__mux2_1
X_05927_ _11221_/Q _06470_/A2 _05925_/X _05926_/X vssd1 vssd1 vccd1 vccd1 _05927_/X
+ sky130_fd_sc_hd__o211a_1
X_09695_ _09673_/B _09672_/Y _09554_/Y vssd1 vssd1 vccd1 vccd1 _09702_/S sky130_fd_sc_hd__o21ai_4
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _08816_/A _08646_/B vssd1 vssd1 vccd1 vccd1 _11179_/D sky130_fd_sc_hd__or2_1
X_05858_ _11153_/Q _06221_/A2 _05856_/X _05857_/X vssd1 vssd1 vccd1 vccd1 _05858_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _11144_/Q _08469_/A _08577_/S vssd1 vssd1 vccd1 vccd1 _08578_/B sky130_fd_sc_hd__mux2_1
X_05789_ _08243_/A _08243_/B vssd1 vssd1 vccd1 vccd1 _05789_/Y sky130_fd_sc_hd__nor2_8
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07528_ _07934_/A _07528_/B vssd1 vssd1 vccd1 vccd1 _10548_/D sky130_fd_sc_hd__or2_1
XFILLER_70_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07459_ _07451_/B _07754_/B _07458_/X vssd1 vssd1 vccd1 vccd1 _10506_/D sky130_fd_sc_hd__a21o_1
XFILLER_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10470_ _11641_/CLK _10470_/D vssd1 vssd1 vccd1 vccd1 _10470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09129_ _09129_/A1 _09127_/B _09129_/B1 vssd1 vssd1 vccd1 vccd1 _09129_/X sky130_fd_sc_hd__a21o_1
XFILLER_109_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11022_ _11733_/CLK _11022_/D vssd1 vssd1 vccd1 vccd1 _11022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ _11457_/CLK _10806_/D vssd1 vssd1 vccd1 vccd1 _10806_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11786_ _11791_/CLK _11786_/D vssd1 vssd1 vccd1 vccd1 _11786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10737_ _11711_/CLK _10737_/D vssd1 vssd1 vccd1 vccd1 _10737_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10668_ _11457_/CLK _10668_/D vssd1 vssd1 vccd1 vccd1 _10668_/Q sky130_fd_sc_hd__dfxtp_1
X_10599_ _11780_/CLK _10599_/D vssd1 vssd1 vccd1 vccd1 _10599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput129 _11609_/Q vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_4
XFILLER_127_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06830_ _10495_/Q _06872_/A2 _06829_/X _06849_/C1 vssd1 vssd1 vccd1 vccd1 _06830_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06761_ _10392_/Q _06860_/A2 _06757_/X _06760_/X vssd1 vssd1 vccd1 vccd1 _06761_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05712_ _11052_/Q _05518_/Y _05524_/Y _11043_/Q vssd1 vssd1 vccd1 vccd1 _05712_/X
+ sky130_fd_sc_hd__a22o_1
X_08500_ _07107_/A _08497_/S _08499_/X _08588_/C1 vssd1 vssd1 vccd1 vccd1 _11100_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06692_ _10759_/Q _07854_/A _07153_/A _11470_/Q _06691_/X vssd1 vssd1 vccd1 vccd1
+ _06692_/X sky130_fd_sc_hd__o221a_1
X_09480_ _09554_/A _09416_/B _09479_/X _09678_/A vssd1 vssd1 vccd1 vccd1 _11603_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08431_ _11056_/Q _08425_/Y _08426_/Y _07013_/X vssd1 vssd1 vccd1 vccd1 _11056_/D
+ sky130_fd_sc_hd__o22a_1
X_05643_ _05643_/A _05643_/B _05643_/C vssd1 vssd1 vccd1 vccd1 _05644_/C sky130_fd_sc_hd__or3_1
XFILLER_24_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08362_ _11024_/Q _08362_/B vssd1 vssd1 vccd1 vccd1 _08362_/X sky130_fd_sc_hd__or2_1
X_05574_ _05628_/A2 _11366_/Q _11363_/Q _05628_/B1 vssd1 vssd1 vccd1 vccd1 _05574_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07313_ _10423_/Q _07301_/Y _07306_/Y _09232_/B2 vssd1 vssd1 vccd1 vccd1 _10423_/D
+ sky130_fd_sc_hd__a22o_1
X_08293_ _10979_/Q _07093_/X _08298_/S vssd1 vssd1 vccd1 vccd1 _10979_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07244_ _07243_/X _10390_/Q _07249_/S vssd1 vssd1 vccd1 vccd1 _10390_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07175_ _07211_/A _09243_/C _07174_/X _07902_/C1 vssd1 vssd1 vccd1 vccd1 _10348_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06126_ _11212_/Q _06126_/B vssd1 vssd1 vccd1 vccd1 _06126_/X sky130_fd_sc_hd__or2_1
XFILLER_30_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06057_ _10439_/Q _06634_/B1 _06731_/B1 _11073_/Q _06550_/C1 vssd1 vssd1 vccd1 vccd1
+ _06057_/X sky130_fd_sc_hd__o221a_2
XFILLER_114_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout301 _08027_/S vssd1 vssd1 vccd1 vccd1 _08035_/S sky130_fd_sc_hd__buf_6
Xfanout312 _07533_/S vssd1 vssd1 vccd1 vccd1 _07513_/S sky130_fd_sc_hd__buf_6
Xfanout323 _07222_/Y vssd1 vssd1 vccd1 vccd1 _07663_/S sky130_fd_sc_hd__buf_8
XFILLER_99_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout334 _07150_/A2 vssd1 vssd1 vccd1 vccd1 _07145_/B sky130_fd_sc_hd__buf_4
XFILLER_8_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout345 _07151_/Y vssd1 vssd1 vccd1 vccd1 _07904_/B sky130_fd_sc_hd__buf_8
Xfanout356 _06997_/Y vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__buf_6
XFILLER_86_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09816_ _09811_/X _09815_/X _08951_/X vssd1 vssd1 vccd1 vccd1 _09824_/S sky130_fd_sc_hd__o21ba_4
Xfanout367 _07232_/B vssd1 vssd1 vccd1 vccd1 _08811_/B2 sky130_fd_sc_hd__buf_6
XFILLER_47_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout378 _07011_/Y vssd1 vssd1 vccd1 vccd1 _08322_/A sky130_fd_sc_hd__buf_12
Xfanout389 _07617_/A vssd1 vssd1 vccd1 vccd1 _07333_/A sky130_fd_sc_hd__buf_6
XFILLER_41_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09747_ _10502_/Q _09879_/A2 _09878_/A2 _10548_/Q vssd1 vssd1 vccd1 vccd1 _09747_/X
+ sky130_fd_sc_hd__a22o_1
X_06959_ _10219_/Q _06958_/X _09416_/A vssd1 vssd1 vccd1 vccd1 _10219_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _09678_/A _09678_/B vssd1 vssd1 vccd1 vccd1 _11634_/D sky130_fd_sc_hd__and2_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08629_ _11169_/Q _08633_/B vssd1 vssd1 vccd1 vccd1 _08629_/X sky130_fd_sc_hd__or2_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ _11641_/CLK _11640_/D vssd1 vssd1 vccd1 vccd1 _11640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11571_ _11573_/CLK _11571_/D vssd1 vssd1 vccd1 vccd1 _11571_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_64_wb_clk_i clkbuf_leaf_69_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11684_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10522_ _10735_/CLK _10522_/D vssd1 vssd1 vccd1 vccd1 _10522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10453_ _11776_/CLK _10453_/D vssd1 vssd1 vccd1 vccd1 _10453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10384_ _10981_/CLK _10384_/D vssd1 vssd1 vccd1 vccd1 _10384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11005_ _11005_/CLK _11005_/D vssd1 vssd1 vccd1 vccd1 _11005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout890 _06194_/A2 vssd1 vssd1 vccd1 vccd1 _06799_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_20_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11769_ _11779_/CLK _11769_/D vssd1 vssd1 vccd1 vccd1 _11769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05290_ _05290_/A _05290_/B _05290_/C _05290_/D vssd1 vssd1 vccd1 vccd1 _05291_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_0__f_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_3_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08980_ _11342_/Q _08972_/X _08979_/X vssd1 vssd1 vccd1 vccd1 _11342_/D sky130_fd_sc_hd__a21o_1
XFILLER_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07931_ _10783_/Q _09208_/B vssd1 vssd1 vccd1 vccd1 _07931_/X sky130_fd_sc_hd__or2_1
XFILLER_151_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07862_ _09090_/A1 _07871_/S _07861_/X _07866_/C1 vssd1 vssd1 vccd1 vccd1 _10749_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09601_ _10379_/Q _09566_/A _09565_/B _10626_/Q vssd1 vssd1 vccd1 vccd1 _09601_/X
+ sky130_fd_sc_hd__a22o_1
X_06813_ _10552_/Q _07440_/A vssd1 vssd1 vccd1 vccd1 _06813_/X sky130_fd_sc_hd__or2_1
XFILLER_151_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07793_ _09129_/A1 _10704_/Q _07817_/S vssd1 vssd1 vccd1 vccd1 _07794_/B sky130_fd_sc_hd__mux2_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09532_ _09492_/B _09500_/B _09508_/A _11621_/Q vssd1 vssd1 vccd1 vccd1 _09532_/X
+ sky130_fd_sc_hd__a31o_1
X_06744_ _10372_/Q _07203_/A _06858_/B1 _10517_/Q _06873_/D1 vssd1 vssd1 vccd1 vccd1
+ _06744_/X sky130_fd_sc_hd__o221a_1
XFILLER_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06675_ _10545_/Q _06728_/B1 _06671_/X _06674_/X vssd1 vssd1 vccd1 vccd1 _06675_/X
+ sky130_fd_sc_hd__o211a_2
X_09463_ _05432_/S _09475_/A _09462_/Y _09407_/A vssd1 vssd1 vccd1 vccd1 _11598_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08414_ _08853_/A1 _11048_/Q _08414_/S vssd1 vssd1 vccd1 vccd1 _08415_/B sky130_fd_sc_hd__mux2_1
X_05626_ _11752_/Q _05626_/A2 _05079_/A _11746_/Q _05625_/X vssd1 vssd1 vccd1 vccd1
+ _05627_/B sky130_fd_sc_hd__a221o_4
X_09394_ _10183_/A0 _11560_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _11560_/D sky130_fd_sc_hd__mux2_1
XFILLER_52_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05557_ _09552_/A1 _11347_/Q _11341_/Q _05078_/A vssd1 vssd1 vccd1 vccd1 _05557_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08345_ _09396_/A0 _08360_/S _08344_/X _08345_/C1 vssd1 vssd1 vccd1 vccd1 _11015_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08276_ _08853_/A1 _10970_/Q _08276_/S vssd1 vssd1 vccd1 vccd1 _08277_/B sky130_fd_sc_hd__mux2_1
XFILLER_138_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05488_ _10233_/Q input44/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05488_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07227_ _07617_/A _07227_/B vssd1 vssd1 vccd1 vccd1 _07227_/X sky130_fd_sc_hd__or2_4
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07158_ _10015_/A0 _10340_/Q _07172_/S vssd1 vssd1 vccd1 vccd1 _07159_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06109_ _10479_/Q _06803_/A2 _06108_/X _06997_/A vssd1 vssd1 vccd1 vccd1 _06109_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07089_ _10300_/Q _07088_/X _07109_/S vssd1 vssd1 vccd1 vccd1 _10300_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_111_wb_clk_i clkbuf_4_10__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11439_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11663_/CLK _11623_/D vssd1 vssd1 vccd1 vccd1 _11623_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11554_ _11763_/CLK _11554_/D vssd1 vssd1 vccd1 vccd1 _11554_/Q sky130_fd_sc_hd__dfxtp_1
X_10505_ _10804_/CLK _10505_/D vssd1 vssd1 vccd1 vccd1 _10505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11485_ _11485_/CLK _11485_/D vssd1 vssd1 vccd1 vccd1 _11485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10436_ _11777_/CLK _10436_/D vssd1 vssd1 vccd1 vccd1 _10436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10367_ _10725_/CLK _10367_/D vssd1 vssd1 vccd1 vccd1 _10367_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _11720_/CLK _10298_/D vssd1 vssd1 vccd1 vccd1 _10298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06460_ _10856_/Q _08054_/A _06458_/X _06459_/X vssd1 vssd1 vccd1 vccd1 _06460_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05411_ _05411_/A _05411_/B _05411_/C _05411_/D vssd1 vssd1 vccd1 vccd1 _05412_/B
+ sky130_fd_sc_hd__or4_2
X_06391_ _10827_/Q _07994_/A _07692_/A _10651_/Q _06390_/X vssd1 vssd1 vccd1 vccd1
+ _06391_/X sky130_fd_sc_hd__o221a_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08130_ _10891_/Q _08637_/C vssd1 vssd1 vccd1 vccd1 _08130_/X sky130_fd_sc_hd__or2_1
X_05342_ _11098_/Q _11097_/Q _05430_/S vssd1 vssd1 vccd1 vccd1 _05345_/B sky130_fd_sc_hd__mux2_1
XFILLER_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08061_ _07061_/A _10856_/Q _08427_/B vssd1 vssd1 vccd1 vccd1 _08062_/B sky130_fd_sc_hd__mux2_1
X_05273_ _10811_/Q _10810_/Q _06967_/A vssd1 vssd1 vccd1 vccd1 _05275_/C sky130_fd_sc_hd__mux2_1
XFILLER_135_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07012_ _09540_/A _08757_/A vssd1 vssd1 vccd1 vccd1 _07012_/Y sky130_fd_sc_hd__nand2_8
XFILLER_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08963_ _09539_/A _09444_/A _09668_/A vssd1 vssd1 vccd1 vccd1 _08963_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07914_ _07928_/A _07914_/B vssd1 vssd1 vccd1 vccd1 _10774_/D sky130_fd_sc_hd__or2_1
XFILLER_97_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08894_ _11304_/Q _08894_/B vssd1 vssd1 vccd1 vccd1 _08894_/X sky130_fd_sc_hd__or2_1
XFILLER_25_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07845_ _07108_/X _10740_/Q _07846_/S vssd1 vssd1 vccd1 vccd1 _10740_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07776_ _07076_/A _07776_/A2 _07204_/Y _10696_/Q _09228_/A vssd1 vssd1 vccd1 vccd1
+ _10696_/D sky130_fd_sc_hd__a221o_1
XFILLER_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09515_ _09522_/B _09515_/B _09515_/C vssd1 vssd1 vccd1 vccd1 _09516_/A sky130_fd_sc_hd__and3_1
X_06727_ _10410_/Q _06727_/B vssd1 vssd1 vccd1 vccd1 _06727_/X sky130_fd_sc_hd__or2_1
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09446_ input21/X input41/X input18/X input27/X _11576_/Q _11577_/Q vssd1 vssd1 vccd1
+ vccd1 _09446_/X sky130_fd_sc_hd__mux4_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06658_ _11204_/Q _10158_/A _09292_/A _11254_/Q vssd1 vssd1 vccd1 vccd1 _06658_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05609_ _05609_/A _05609_/B vssd1 vssd1 vccd1 vccd1 _05609_/Y sky130_fd_sc_hd__nor2_8
XFILLER_12_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09377_ _09995_/A1 _09359_/X _09376_/X _09995_/C1 vssd1 vssd1 vccd1 vccd1 _11546_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06589_ _11101_/Q _06589_/A2 _06588_/X _07690_/B vssd1 vssd1 vccd1 vccd1 _06589_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08328_ _11003_/Q _08322_/Y _08325_/Y _07229_/X vssd1 vssd1 vccd1 vccd1 _11003_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08259_ _08875_/A _08259_/B vssd1 vssd1 vccd1 vccd1 _10961_/D sky130_fd_sc_hd__or2_1
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ _11270_/CLK _11270_/D vssd1 vssd1 vccd1 vccd1 _11270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10221_ _11573_/CLK _10221_/D vssd1 vssd1 vccd1 vccd1 _10221_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_134_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10152_ _11789_/Q _10154_/B vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__or2_1
XFILLER_133_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10083_ _11743_/Q _07227_/X _10085_/S vssd1 vssd1 vccd1 vccd1 _11743_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10985_ _11633_/CLK _10985_/D vssd1 vssd1 vccd1 vccd1 _10985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11606_ _11675_/CLK _11606_/D vssd1 vssd1 vccd1 vccd1 _11606_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11537_ _11733_/CLK _11537_/D vssd1 vssd1 vccd1 vccd1 _11537_/Q sky130_fd_sc_hd__dfxtp_1
X_11468_ _11474_/CLK _11468_/D vssd1 vssd1 vccd1 vccd1 _11468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10419_ _11233_/CLK _10419_/D vssd1 vssd1 vccd1 vccd1 _10419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11399_ _11462_/CLK _11399_/D vssd1 vssd1 vccd1 vccd1 _11399_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05960_ _11425_/Q _08668_/A _05959_/X _06670_/D1 vssd1 vssd1 vccd1 vccd1 _05960_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05891_ _11678_/Q _09977_/A _05887_/X _05890_/X vssd1 vssd1 vccd1 vccd1 _05891_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07630_ _08810_/A _07630_/B vssd1 vssd1 vccd1 vccd1 _07630_/Y sky130_fd_sc_hd__nor2_2
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07561_ _08876_/A0 _10564_/Q _07589_/S vssd1 vssd1 vccd1 vccd1 _07562_/B sky130_fd_sc_hd__mux2_1
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09300_ _09985_/A1 _09310_/B _10166_/B1 vssd1 vssd1 vccd1 vccd1 _09300_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06512_ _10921_/Q _06591_/A2 _06126_/B _11217_/Q _06511_/X vssd1 vssd1 vccd1 vccd1
+ _06512_/X sky130_fd_sc_hd__o221a_1
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07492_ _07248_/X _10528_/Q _07496_/S vssd1 vssd1 vccd1 vccd1 _10528_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09231_ _11465_/Q _09226_/Y _09229_/Y _07016_/X vssd1 vssd1 vccd1 vccd1 _11465_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06443_ _11043_/Q _09059_/A _08971_/A _10965_/Q vssd1 vssd1 vccd1 vccd1 _06443_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09162_ _11425_/Q _09154_/X _09161_/X vssd1 vssd1 vccd1 vccd1 _11425_/D sky130_fd_sc_hd__a21o_1
X_06374_ _06374_/A _06374_/B _06374_/C vssd1 vssd1 vccd1 vccd1 _06374_/X sky130_fd_sc_hd__and3_4
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08113_ _10882_/Q _08120_/S _07642_/S _07098_/B vssd1 vssd1 vccd1 vccd1 _10882_/D
+ sky130_fd_sc_hd__o22a_1
X_05325_ _10461_/Q _10848_/Q _05385_/S vssd1 vssd1 vccd1 vccd1 _05329_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09093_ _09283_/A1 _09099_/B _08873_/A vssd1 vssd1 vccd1 vccd1 _09093_/X sky130_fd_sc_hd__a21o_1
X_08044_ _10847_/Q _08051_/S _07365_/Y _07098_/B vssd1 vssd1 vccd1 vccd1 _10847_/D
+ sky130_fd_sc_hd__o22a_1
X_05256_ _10978_/Q _10977_/Q _05429_/S vssd1 vssd1 vccd1 vccd1 _05258_/C sky130_fd_sc_hd__mux2_1
XFILLER_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05187_ _10843_/Q _10842_/Q _05471_/A vssd1 vssd1 vccd1 vccd1 _05189_/C sky130_fd_sc_hd__mux2_1
XFILLER_131_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09995_ _09995_/A1 _09977_/X _09994_/X _09995_/C1 vssd1 vssd1 vccd1 vccd1 _11684_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08946_ _11332_/Q _08946_/B vssd1 vssd1 vccd1 vccd1 _08946_/X sky130_fd_sc_hd__or2_1
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08877_ _08941_/A _08877_/B vssd1 vssd1 vccd1 vccd1 _11295_/D sky130_fd_sc_hd__or2_1
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07828_ _07059_/A _07839_/A2 _07821_/A _10723_/Q vssd1 vssd1 vccd1 vccd1 _10723_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07759_ _07039_/A _07761_/A2 _07758_/X _09201_/A1 vssd1 vssd1 vccd1 vccd1 _10680_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10770_ _10805_/CLK _10770_/D vssd1 vssd1 vccd1 vccd1 _10770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09429_ _09540_/A _09428_/X _09703_/A vssd1 vssd1 vccd1 vccd1 _11587_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11322_ _11332_/CLK _11322_/D vssd1 vssd1 vccd1 vccd1 _11322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11253_ _11329_/CLK _11253_/D vssd1 vssd1 vccd1 vccd1 _11253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10204_ _11758_/CLK _10204_/D vssd1 vssd1 vccd1 vccd1 _10204_/Q sky130_fd_sc_hd__dfxtp_1
X_11184_ _11224_/CLK _11184_/D vssd1 vssd1 vccd1 vccd1 _11184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10135_ _10135_/A0 _11781_/Q _10135_/S vssd1 vssd1 vccd1 vccd1 _11781_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10066_ _10113_/A0 _11727_/Q _10071_/S vssd1 vssd1 vccd1 vccd1 _11727_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10968_ _11243_/CLK _10968_/D vssd1 vssd1 vccd1 vccd1 _10968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10899_ _11601_/CLK _10899_/D vssd1 vssd1 vccd1 vccd1 _10899_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05110_ _10606_/Q _10605_/Q _05398_/S vssd1 vssd1 vccd1 vccd1 _05112_/C sky130_fd_sc_hd__mux2_1
XFILLER_156_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06090_ _11374_/Q _09038_/A _09110_/A _11407_/Q _06089_/X vssd1 vssd1 vccd1 vccd1
+ _06090_/X sky130_fd_sc_hd__o221a_1
XFILLER_8_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout708 _07297_/Y vssd1 vssd1 vccd1 vccd1 _10136_/C sky130_fd_sc_hd__buf_6
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout719 fanout726/X vssd1 vssd1 vccd1 vccd1 _06105_/B1 sky130_fd_sc_hd__buf_4
XFILLER_98_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _11256_/Q _08804_/B vssd1 vssd1 vccd1 vccd1 _08800_/X sky130_fd_sc_hd__or2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09780_ _11648_/Q _09771_/Y _09779_/X _09554_/B _09406_/B vssd1 vssd1 vccd1 vccd1
+ _09780_/X sky130_fd_sc_hd__o221a_1
X_06992_ _10263_/Q _06976_/X _06991_/X vssd1 vssd1 vccd1 vccd1 _10263_/D sky130_fd_sc_hd__a21o_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _07010_/A _08748_/S _08730_/X _08821_/A vssd1 vssd1 vccd1 vccd1 _11222_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05943_ _11145_/Q _07692_/A _05941_/X _05942_/X vssd1 vssd1 vccd1 vccd1 _05943_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08662_ _11186_/Q _08663_/S _08661_/X _08662_/C1 vssd1 vssd1 vccd1 vccd1 _11186_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05874_ _10634_/Q _06453_/B1 _05873_/X _06265_/C1 vssd1 vssd1 vccd1 vccd1 _05874_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07613_ _07613_/A _08037_/B vssd1 vssd1 vccd1 vccd1 _07613_/Y sky130_fd_sc_hd__nor2_2
XFILLER_148_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08593_ _09038_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08633_/B sky130_fd_sc_hd__nor2_8
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07544_ _08536_/A _07544_/B vssd1 vssd1 vccd1 vccd1 _10555_/D sky130_fd_sc_hd__or2_1
XFILLER_22_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07475_ _07070_/A _10516_/Q _07477_/S vssd1 vssd1 vccd1 vccd1 _07476_/B sky130_fd_sc_hd__mux2_1
X_09214_ _09214_/A _09214_/B _09221_/C vssd1 vssd1 vccd1 vccd1 _09214_/X sky130_fd_sc_hd__or3_1
X_06426_ _11309_/Q _06640_/B1 _08469_/B _10983_/Q vssd1 vssd1 vccd1 vccd1 _06426_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_50_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09145_ _11418_/Q _09149_/B vssd1 vssd1 vccd1 vccd1 _09145_/X sky130_fd_sc_hd__or2_1
X_06357_ _11378_/Q _09038_/A _06356_/X _06357_/C1 vssd1 vssd1 vccd1 vccd1 _06357_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05308_ _11012_/Q _11011_/Q _11594_/Q vssd1 vssd1 vccd1 vccd1 _05312_/A sky130_fd_sc_hd__mux2_1
X_09076_ _11386_/Q _09060_/X _09075_/X vssd1 vssd1 vccd1 vccd1 _11386_/D sky130_fd_sc_hd__a21o_1
X_06288_ _11871_/A _08243_/B vssd1 vssd1 vccd1 vccd1 _06900_/A sky130_fd_sc_hd__nor2_2
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08027_ _09995_/A1 _10838_/Q _08027_/S vssd1 vssd1 vccd1 vccd1 _08028_/B sky130_fd_sc_hd__mux2_1
X_05239_ _10788_/Q _10862_/Q _06939_/A vssd1 vssd1 vccd1 vccd1 _05239_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_89_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11665_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09978_ _10161_/A1 _09994_/B _08851_/A vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10981_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08929_ _08929_/A1 _08945_/A2 _08928_/X _08947_/C1 vssd1 vssd1 vccd1 vccd1 _11323_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _11871_/A vssd1 vssd1 vccd1 vccd1 _11871_/X sky130_fd_sc_hd__buf_2
XFILLER_79_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10822_ _11633_/CLK _10822_/D vssd1 vssd1 vccd1 vccd1 _10822_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10753_ _10808_/CLK _10753_/D vssd1 vssd1 vccd1 vccd1 _10753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10684_ _11713_/CLK _10684_/D vssd1 vssd1 vccd1 vccd1 _10684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11305_ _11308_/CLK _11305_/D vssd1 vssd1 vccd1 vccd1 _11305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11236_ _11366_/CLK _11236_/D vssd1 vssd1 vccd1 vccd1 _11236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11167_ _11329_/CLK _11167_/D vssd1 vssd1 vccd1 vccd1 _11167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10118_ _10118_/A0 _11765_/Q _10118_/S vssd1 vssd1 vccd1 vccd1 _11765_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11098_ _11607_/CLK _11098_/D vssd1 vssd1 vccd1 vccd1 _11098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10049_ _11716_/Q _07034_/A _10051_/S vssd1 vssd1 vccd1 vccd1 _10050_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05590_ _05626_/A2 _10199_/Q _10194_/Q _05630_/B1 _05589_/X vssd1 vssd1 vccd1 vccd1
+ _05591_/B sky130_fd_sc_hd__a221o_4
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07260_ _07790_/A _07260_/B vssd1 vssd1 vccd1 vccd1 _10398_/D sky130_fd_sc_hd__or2_1
XFILLER_91_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06211_ _06663_/A _10228_/Q _06622_/B2 _06210_/X vssd1 vssd1 vccd1 vccd1 _10228_/D
+ sky130_fd_sc_hd__a31o_1
X_07191_ _07309_/A _07191_/B vssd1 vssd1 vccd1 vccd1 _07192_/A sky130_fd_sc_hd__nor2_8
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06142_ _07151_/B _06115_/X _06120_/X _06104_/X vssd1 vssd1 vccd1 vccd1 _06142_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_144_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06073_ _11147_/Q _06161_/A2 _06071_/X _06072_/X vssd1 vssd1 vccd1 vccd1 _06073_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09901_ _11719_/Q _09571_/A _09909_/A2 _11722_/Q _09900_/X vssd1 vssd1 vccd1 vccd1
+ _09901_/X sky130_fd_sc_hd__a221o_1
XFILLER_132_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout505 _09048_/C1 vssd1 vssd1 vccd1 vccd1 _09122_/C1 sky130_fd_sc_hd__buf_4
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout516 _08050_/A vssd1 vssd1 vccd1 vccd1 _08745_/A sky130_fd_sc_hd__buf_4
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _09831_/X _11657_/Q _09832_/S vssd1 vssd1 vccd1 vccd1 _09833_/B sky130_fd_sc_hd__mux2_1
Xfanout527 _08590_/A vssd1 vssd1 vccd1 vccd1 _08835_/A sky130_fd_sc_hd__buf_4
Xfanout538 _10056_/A vssd1 vssd1 vccd1 vccd1 _10043_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout549 _07790_/A vssd1 vssd1 vccd1 vccd1 _07916_/A sky130_fd_sc_hd__buf_4
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ input7/X _09740_/Y _09762_/X vssd1 vssd1 vccd1 vccd1 _09763_/X sky130_fd_sc_hd__a21o_1
X_06975_ _07939_/A _08649_/B _10158_/B vssd1 vssd1 vccd1 vccd1 _06995_/B sky130_fd_sc_hd__and3_4
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08714_ _11212_/Q _08718_/S _07852_/S _07617_/B vssd1 vssd1 vccd1 vccd1 _11212_/D
+ sky130_fd_sc_hd__o22a_1
X_05926_ _10462_/Q _06642_/A2 _08469_/B _10977_/Q vssd1 vssd1 vccd1 vccd1 _05926_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_67_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09694_ _09703_/A _09694_/B vssd1 vssd1 vccd1 vccd1 _11638_/D sky130_fd_sc_hd__or2_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _11179_/Q _08818_/A1 _08645_/S vssd1 vssd1 vccd1 vccd1 _08646_/B sky130_fd_sc_hd__mux2_1
X_05857_ _11034_/Q _06735_/A2 _06717_/B1 _10956_/Q vssd1 vssd1 vccd1 vccd1 _05857_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08576_ _08749_/A _08576_/B vssd1 vssd1 vccd1 vccd1 _11143_/D sky130_fd_sc_hd__or2_1
XFILLER_39_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05788_ _11189_/Q _06736_/A2 _09038_/A _11152_/Q vssd1 vssd1 vccd1 vccd1 _05788_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07527_ _07034_/A _10548_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _07528_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_136_wb_clk_i clkbuf_4_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11133_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07458_ _10506_/Q _09243_/B _07755_/A2 _09192_/A vssd1 vssd1 vccd1 vccd1 _07458_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06409_ _11609_/Q _06665_/A2 _06406_/X _06853_/A3 _06408_/X vssd1 vssd1 vccd1 vccd1
+ _10231_/D sky130_fd_sc_hd__a221o_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07389_ _08749_/A _07389_/B vssd1 vssd1 vccd1 vccd1 _10470_/D sky130_fd_sc_hd__or2_1
XFILLER_124_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09128_ _09289_/A1 _09110_/X _09127_/X _09289_/C1 vssd1 vssd1 vccd1 vccd1 _11410_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09059_ _09059_/A _10136_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09077_/B sky130_fd_sc_hd__and3_4
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11021_ _11023_/CLK _11021_/D vssd1 vssd1 vccd1 vccd1 _11021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1130 vssd1 vssd1 vccd1 vccd1 io_oeb[7] wrapped_tms1x00_1130/LO sky130_fd_sc_hd__conb_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10805_ _10805_/CLK _10805_/D vssd1 vssd1 vccd1 vccd1 _10805_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11785_ _11809_/CLK _11785_/D vssd1 vssd1 vccd1 vccd1 _11785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10736_ _11745_/CLK _10736_/D vssd1 vssd1 vccd1 vccd1 _10736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ _10782_/CLK _10667_/D vssd1 vssd1 vccd1 vccd1 _10667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10598_ _11766_/CLK _10598_/D vssd1 vssd1 vccd1 vccd1 _10598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11219_ _11779_/CLK _11219_/D vssd1 vssd1 vccd1 vccd1 _11219_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06760_ _10732_/Q _07819_/A _06759_/X _06849_/C1 vssd1 vssd1 vccd1 vccd1 _06760_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05711_ _11051_/Q _05591_/Y _05633_/Y _11034_/Q _05710_/X vssd1 vssd1 vccd1 vccd1
+ _05716_/B sky130_fd_sc_hd__a221o_2
X_06691_ _10780_/Q _06862_/A2 _06877_/B1 _10571_/Q vssd1 vssd1 vccd1 vccd1 _06691_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_149_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08430_ _11055_/Q _08424_/Y _08427_/Y _07008_/X vssd1 vssd1 vccd1 vccd1 _11055_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05642_ _11328_/Q _05561_/Y _05585_/Y _11327_/Q _05641_/X vssd1 vssd1 vccd1 vccd1
+ _05643_/C sky130_fd_sc_hd__a221o_1
X_08361_ _08835_/A _08361_/B vssd1 vssd1 vccd1 vccd1 _11023_/D sky130_fd_sc_hd__or2_1
X_05573_ _05573_/A _05573_/B vssd1 vssd1 vccd1 vccd1 _05573_/Y sky130_fd_sc_hd__nor2_8
X_07312_ _10422_/Q _07302_/Y _07305_/Y _07232_/X vssd1 vssd1 vccd1 vccd1 _10422_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ _10978_/Q _07227_/X _08298_/S vssd1 vssd1 vccd1 vccd1 _10978_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07243_ _09206_/A _07243_/B vssd1 vssd1 vccd1 vccd1 _07243_/X sky130_fd_sc_hd__and2_1
XFILLER_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07174_ _10348_/Q _09228_/B vssd1 vssd1 vccd1 vccd1 _07174_/X sky130_fd_sc_hd__or2_1
XFILLER_145_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06125_ _06125_/A _06125_/B _06125_/C vssd1 vssd1 vccd1 vccd1 _06125_/X sky130_fd_sc_hd__and3_1
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06056_ _10913_/Q _06591_/A2 _06637_/A2 _11211_/Q _06055_/X vssd1 vssd1 vccd1 vccd1
+ _06059_/A sky130_fd_sc_hd__o221a_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout302 _07557_/S vssd1 vssd1 vccd1 vccd1 _07591_/S sky130_fd_sc_hd__buf_8
XFILLER_87_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout313 _07535_/S vssd1 vssd1 vccd1 vccd1 _07533_/S sky130_fd_sc_hd__buf_6
Xfanout324 _07222_/Y vssd1 vssd1 vccd1 vccd1 _07665_/S sky130_fd_sc_hd__buf_6
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout335 _07110_/Y vssd1 vssd1 vccd1 vccd1 _07150_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_28_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout346 _07151_/Y vssd1 vssd1 vccd1 vccd1 _07854_/B sky130_fd_sc_hd__buf_6
Xfanout357 _09271_/B vssd1 vssd1 vccd1 vccd1 _10137_/B sky130_fd_sc_hd__buf_6
X_09815_ _09815_/A _09815_/B _09815_/C _09815_/D vssd1 vssd1 vccd1 vccd1 _09815_/X
+ sky130_fd_sc_hd__or4_1
Xfanout368 _07018_/X vssd1 vssd1 vccd1 vccd1 _07232_/B sky130_fd_sc_hd__buf_8
XFILLER_86_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout379 _09214_/B vssd1 vssd1 vccd1 vccd1 _07441_/A sky130_fd_sc_hd__buf_6
XFILLER_46_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09746_ _10547_/Q _09879_/B1 _09878_/B1 _10500_/Q _09745_/X vssd1 vssd1 vccd1 vccd1
+ _09749_/C sky130_fd_sc_hd__a221o_1
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06958_ _11663_/Q _05474_/B _06955_/X _05474_/A _06957_/X vssd1 vssd1 vccd1 vccd1
+ _06958_/X sky130_fd_sc_hd__a221o_4
XFILLER_132_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05909_ _10267_/Q _06999_/A _06857_/B1 _11698_/Q vssd1 vssd1 vccd1 vccd1 _05909_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09540_/A _09554_/Y _09675_/X _09676_/Y _11634_/Q vssd1 vssd1 vccd1 vccd1
+ _09678_/B sky130_fd_sc_hd__a32o_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06889_ _07048_/A _08970_/S _06884_/Y _10213_/Q vssd1 vssd1 vccd1 vccd1 _10213_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _09216_/A0 _08623_/S _08627_/X _08921_/C1 vssd1 vssd1 vccd1 vccd1 _11168_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _08821_/A _08559_/B vssd1 vssd1 vccd1 vccd1 _11134_/D sky130_fd_sc_hd__and2_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11570_ _11573_/CLK _11570_/D vssd1 vssd1 vccd1 vccd1 _11570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10521_ _11713_/CLK _10521_/D vssd1 vssd1 vccd1 vccd1 _10521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10452_ _11310_/CLK _10452_/D vssd1 vssd1 vccd1 vccd1 _10452_/Q sky130_fd_sc_hd__dfxtp_1
X_10383_ _11661_/CLK _10383_/D vssd1 vssd1 vccd1 vccd1 _10383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11756_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ _11234_/CLK _11004_/D vssd1 vssd1 vccd1 vccd1 _11004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout880 _06370_/A2 vssd1 vssd1 vccd1 vccd1 _07202_/A sky130_fd_sc_hd__buf_6
Xfanout891 _06862_/A2 vssd1 vssd1 vccd1 vccd1 _06875_/A2 sky130_fd_sc_hd__buf_6
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11768_ _11768_/CLK _11768_/D vssd1 vssd1 vccd1 vccd1 _11768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10719_ _11706_/CLK _10719_/D vssd1 vssd1 vccd1 vccd1 _10719_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11699_ _11702_/CLK _11699_/D vssd1 vssd1 vccd1 vccd1 _11699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ _07930_/A _07930_/B vssd1 vssd1 vccd1 vccd1 _10782_/D sky130_fd_sc_hd__or2_1
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07861_ _10749_/Q _07883_/B vssd1 vssd1 vccd1 vccd1 _07861_/X sky130_fd_sc_hd__or2_1
XFILLER_84_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09600_ _09600_/A _09600_/B vssd1 vssd1 vccd1 vccd1 _09600_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06812_ _11631_/Q _06704_/B _06811_/X vssd1 vssd1 vccd1 vccd1 _10246_/D sky130_fd_sc_hd__a21o_1
XFILLER_68_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07792_ _07926_/A _07792_/B vssd1 vssd1 vccd1 vccd1 _10703_/D sky130_fd_sc_hd__or2_1
X_09531_ _09525_/A _09528_/B _09504_/Y _09530_/X _09825_/A vssd1 vssd1 vccd1 vccd1
+ _11620_/D sky130_fd_sc_hd__o311a_1
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06743_ _06743_/A _06743_/B vssd1 vssd1 vccd1 vccd1 _06743_/X sky130_fd_sc_hd__and2_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09462_ _09475_/A _09462_/B vssd1 vssd1 vccd1 vccd1 _09462_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06674_ _10669_/Q _06674_/A2 _06673_/X _06808_/C1 vssd1 vssd1 vccd1 vccd1 _06674_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ _08684_/A _08413_/B vssd1 vssd1 vccd1 vccd1 _11047_/D sky130_fd_sc_hd__or2_1
X_05625_ _11755_/Q _05631_/A2 _05631_/B1 _11751_/Q _05623_/X vssd1 vssd1 vccd1 vccd1
+ _05625_/X sky130_fd_sc_hd__a221o_1
X_09393_ _09393_/A0 _11559_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _11559_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08344_ _11015_/Q _08362_/B vssd1 vssd1 vccd1 vccd1 _08344_/X sky130_fd_sc_hd__or2_1
X_05556_ _05616_/A1 _11346_/Q _11343_/Q _05077_/A vssd1 vssd1 vccd1 vccd1 _05556_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08275_ _08536_/A _08275_/B vssd1 vssd1 vccd1 vccd1 _10969_/D sky130_fd_sc_hd__or2_1
X_05487_ _10232_/Q input43/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05487_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07226_ _08441_/B2 _10380_/Q _07246_/S vssd1 vssd1 vccd1 vccd1 _10380_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07157_ _07928_/A _07157_/B vssd1 vssd1 vccd1 vccd1 _10339_/D sky130_fd_sc_hd__or2_1
XFILLER_69_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06108_ _10509_/Q _06999_/A _07539_/A _10315_/Q _06107_/X vssd1 vssd1 vccd1 vccd1
+ _06108_/X sky130_fd_sc_hd__o221a_1
XFILLER_65_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07088_ _07318_/A _07324_/B vssd1 vssd1 vccd1 vccd1 _07088_/X sky130_fd_sc_hd__or2_4
XFILLER_65_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06039_ _07690_/A _06033_/X _06038_/X _08243_/A _06028_/X vssd1 vssd1 vccd1 vccd1
+ _06039_/X sky130_fd_sc_hd__o311a_2
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09729_ _10339_/Q _09875_/B1 _09878_/B1 _11470_/Q vssd1 vssd1 vccd1 vccd1 _09729_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11622_ _11622_/CLK _11622_/D vssd1 vssd1 vccd1 vccd1 _11622_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ _11763_/CLK _11553_/D vssd1 vssd1 vccd1 vccd1 _11553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10504_ _11450_/CLK _10504_/D vssd1 vssd1 vccd1 vccd1 _10504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11484_ _11809_/CLK _11484_/D vssd1 vssd1 vccd1 vccd1 _11484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10435_ _11766_/CLK _10435_/D vssd1 vssd1 vccd1 vccd1 _10435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10366_ _11698_/CLK _10366_/D vssd1 vssd1 vccd1 vccd1 _10366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10297_ _11698_/CLK _10297_/D vssd1 vssd1 vccd1 vccd1 _10297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05410_ _10588_/Q _10587_/Q _06945_/B vssd1 vssd1 vccd1 vccd1 _05411_/D sky130_fd_sc_hd__mux2_1
X_06390_ _10854_/Q _06631_/A2 _06628_/B1 _11272_/Q vssd1 vssd1 vccd1 vccd1 _06390_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05341_ _11090_/Q _11089_/Q _06939_/A vssd1 vssd1 vccd1 vccd1 _05345_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08060_ _07059_/A _08427_/B _08059_/X _08831_/C1 vssd1 vssd1 vccd1 vccd1 _10855_/D
+ sky130_fd_sc_hd__o211a_1
X_05272_ _10815_/Q _10814_/Q _05392_/S vssd1 vssd1 vccd1 vccd1 _05275_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07011_ _09668_/A _07011_/B vssd1 vssd1 vccd1 vccd1 _07011_/Y sky130_fd_sc_hd__nor2_4
XFILLER_31_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08962_ _11333_/Q _08965_/A _08961_/Y _09833_/A vssd1 vssd1 vccd1 vccd1 _11333_/D
+ sky130_fd_sc_hd__o211a_1
X_07913_ _08929_/A1 _10774_/Q _09221_/C vssd1 vssd1 vccd1 vccd1 _07914_/B sky130_fd_sc_hd__mux2_1
XFILLER_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08893_ _08893_/A1 _08884_/S _08892_/X _09092_/C1 vssd1 vssd1 vccd1 vccd1 _11303_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07844_ _07316_/X _10739_/Q _07846_/S vssd1 vssd1 vccd1 vccd1 _10739_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07775_ _07141_/X _07776_/A2 _07204_/Y _10695_/Q _09214_/B vssd1 vssd1 vccd1 vccd1
+ _10695_/D sky130_fd_sc_hd__a221o_1
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09514_ _09492_/B _09502_/B _09512_/Y _09513_/X _09529_/A vssd1 vssd1 vccd1 vccd1
+ _11614_/D sky130_fd_sc_hd__o311a_1
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06726_ _10349_/Q _07153_/A vssd1 vssd1 vccd1 vccd1 _06726_/X sky130_fd_sc_hd__or2_1
X_09445_ _09407_/B _09443_/X _09444_/Y _09414_/S vssd1 vssd1 vccd1 vccd1 _11594_/D
+ sky130_fd_sc_hd__a22o_1
X_06657_ _11328_/Q _10086_/A _10136_/A _11300_/Q _08243_/B vssd1 vssd1 vccd1 vccd1
+ _06657_/X sky130_fd_sc_hd__a221o_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05608_ _05626_/A2 _11544_/Q _11539_/Q _05630_/B1 _05607_/X vssd1 vssd1 vccd1 vccd1
+ _05609_/B sky130_fd_sc_hd__a221o_4
X_09376_ _11546_/Q _09376_/B vssd1 vssd1 vccd1 vccd1 _09376_/X sky130_fd_sc_hd__or2_1
XFILLER_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06588_ _10947_/Q _06630_/A2 _06632_/A2 _10899_/Q _06587_/X vssd1 vssd1 vccd1 vccd1
+ _06588_/X sky130_fd_sc_hd__o221a_2
XFILLER_21_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08327_ _11002_/Q _08322_/Y _08325_/Y _07008_/X vssd1 vssd1 vccd1 vccd1 _11002_/D
+ sky130_fd_sc_hd__a22o_1
X_05539_ _05629_/A2 _11357_/Q _11351_/Q _05629_/B1 vssd1 vssd1 vccd1 vccd1 _05539_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_138_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08258_ _09124_/A1 _10961_/Q _08276_/S vssd1 vssd1 vccd1 vccd1 _08259_/B sky130_fd_sc_hd__mux2_1
XFILLER_138_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07209_ _07061_/A _07205_/B _07773_/S _10367_/Q vssd1 vssd1 vccd1 vccd1 _10367_/D
+ sky130_fd_sc_hd__o22a_1
X_08189_ _10929_/Q _10128_/A0 _08197_/S vssd1 vssd1 vccd1 vccd1 _08190_/B sky130_fd_sc_hd__mux2_1
XFILLER_134_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10220_ _11573_/CLK _10220_/D vssd1 vssd1 vccd1 vccd1 _10220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10151_ _11788_/Q _10137_/X _10150_/X vssd1 vssd1 vccd1 vccd1 _11788_/D sky130_fd_sc_hd__a21o_1
XFILLER_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10082_ _10118_/A0 _11742_/Q _10082_/S vssd1 vssd1 vccd1 vccd1 _11742_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10984_ _11310_/CLK _10984_/D vssd1 vssd1 vccd1 vccd1 _10984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11605_ _11675_/CLK _11605_/D vssd1 vssd1 vccd1 vccd1 _11605_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11536_ _11765_/CLK _11536_/D vssd1 vssd1 vccd1 vccd1 _11536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11467_ _11471_/CLK _11467_/D vssd1 vssd1 vccd1 vccd1 _11467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10418_ _11233_/CLK _10418_/D vssd1 vssd1 vccd1 vccd1 _10418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11398_ _11410_/CLK _11398_/D vssd1 vssd1 vccd1 vccd1 _11398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _10785_/CLK _10349_/D vssd1 vssd1 vccd1 vccd1 _10349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05890_ _11540_/Q _09359_/A _05888_/X _05889_/X vssd1 vssd1 vccd1 vccd1 _05890_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ _08781_/A _07560_/B vssd1 vssd1 vccd1 vccd1 _10563_/D sky130_fd_sc_hd__or2_1
XFILLER_59_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06511_ _11133_/Q _07222_/A _07819_/A _10308_/Q vssd1 vssd1 vccd1 vccd1 _06511_/X
+ sky130_fd_sc_hd__o22a_2
X_07491_ _07026_/X _10527_/Q _07491_/S vssd1 vssd1 vccd1 vccd1 _10527_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09230_ _11464_/Q _09226_/Y _09229_/Y _07617_/X vssd1 vssd1 vccd1 vccd1 _11464_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06442_ _06436_/X _06441_/X _11872_/A vssd1 vssd1 vccd1 vccd1 _06442_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ _09985_/A1 _09171_/B _08771_/A vssd1 vssd1 vccd1 vccd1 _09161_/X sky130_fd_sc_hd__a21o_1
X_06373_ _10287_/Q _07046_/A _06373_/B1 _10318_/Q _06370_/X vssd1 vssd1 vccd1 vccd1
+ _06374_/C sky130_fd_sc_hd__o221a_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08112_ _08193_/A _08112_/B vssd1 vssd1 vccd1 vccd1 _10881_/D sky130_fd_sc_hd__or2_1
X_05324_ _05324_/A _05324_/B vssd1 vssd1 vccd1 vccd1 _05324_/Y sky130_fd_sc_hd__nor2_8
X_09092_ _09280_/A1 _09082_/X _09091_/X _09092_/C1 vssd1 vssd1 vccd1 vccd1 _11393_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08043_ _08196_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _10846_/D sky130_fd_sc_hd__or2_1
XFILLER_107_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05255_ _11084_/Q _11083_/Q _05397_/S vssd1 vssd1 vccd1 vccd1 _05258_/B sky130_fd_sc_hd__mux2_1
XFILLER_134_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05186_ _10596_/Q _10595_/Q _05419_/S vssd1 vssd1 vccd1 vccd1 _05189_/B sky130_fd_sc_hd__mux2_1
XFILLER_1_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09994_ _11684_/Q _09994_/B vssd1 vssd1 vccd1 vccd1 _09994_/X sky130_fd_sc_hd__or2_1
XFILLER_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08945_ input97/X _08945_/A2 _08944_/X _09122_/C1 vssd1 vssd1 vccd1 vccd1 _11331_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08876_ _08876_/A0 _11295_/Q _08890_/S vssd1 vssd1 vccd1 vccd1 _08877_/B sky130_fd_sc_hd__mux2_1
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07827_ _07057_/A _07827_/A2 _10010_/B _07821_/Y _10722_/Q vssd1 vssd1 vccd1 vccd1
+ _10722_/D sky130_fd_sc_hd__o32a_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07758_ _10680_/Q _07760_/B vssd1 vssd1 vccd1 vccd1 _07758_/X sky130_fd_sc_hd__or2_1
XFILLER_38_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06709_ _11471_/Q _07153_/A _06705_/X _06708_/X vssd1 vssd1 vccd1 vccd1 _06709_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07689_ _07689_/A _07689_/B vssd1 vssd1 vccd1 vccd1 _07689_/Y sky130_fd_sc_hd__nor2_8
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09428_ input1/X _10217_/Q _10213_/Q vssd1 vssd1 vccd1 vccd1 _09428_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09359_ _09359_/A _10137_/B _10159_/C vssd1 vssd1 vccd1 vccd1 _09359_/X sky130_fd_sc_hd__or3_4
XFILLER_139_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11321_ _11393_/CLK _11321_/D vssd1 vssd1 vccd1 vccd1 _11321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11252_ _11812_/CLK _11252_/D vssd1 vssd1 vccd1 vccd1 _11252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10203_ _11809_/CLK _10203_/D vssd1 vssd1 vccd1 vccd1 _10203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11183_ _11629_/CLK _11183_/D vssd1 vssd1 vccd1 vccd1 _11183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ _10134_/A0 _11780_/Q _10134_/S vssd1 vssd1 vccd1 vccd1 _11780_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10065_ _10112_/A0 _11726_/Q _10071_/S vssd1 vssd1 vccd1 vccd1 _11726_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10967_ _11243_/CLK _10967_/D vssd1 vssd1 vccd1 vccd1 _10967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10898_ _11604_/CLK _10898_/D vssd1 vssd1 vccd1 vccd1 _10898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11519_ _11685_/CLK _11519_/D vssd1 vssd1 vccd1 vccd1 _11519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout709 _07297_/Y vssd1 vssd1 vccd1 vccd1 _10158_/C sky130_fd_sc_hd__clkbuf_4
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _10153_/A1 _06995_/B _08664_/A vssd1 vssd1 vccd1 vccd1 _06991_/X sky130_fd_sc_hd__a21o_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _11222_/Q _08750_/B vssd1 vssd1 vccd1 vccd1 _08730_/X sky130_fd_sc_hd__or2_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05942_ _10937_/Q _10061_/A _06459_/B1 _11013_/Q vssd1 vssd1 vccd1 vccd1 _05942_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_112_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08661_ _08661_/A _09249_/A _10119_/B _10087_/C vssd1 vssd1 vccd1 vccd1 _08661_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_61_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05873_ _10582_/Q _06454_/A2 _06455_/B1 _10901_/Q _05872_/X vssd1 vssd1 vccd1 vccd1
+ _05873_/X sky130_fd_sc_hd__o221a_2
XFILLER_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07612_ _09977_/A _08230_/B _10159_/C vssd1 vssd1 vccd1 vccd1 _08027_/S sky130_fd_sc_hd__or3_4
X_08592_ _08665_/A _08589_/S _08591_/X _08662_/C1 vssd1 vssd1 vccd1 vccd1 _11151_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07543_ _10013_/A0 _10555_/Q _07591_/S vssd1 vssd1 vccd1 vccd1 _07544_/B sky130_fd_sc_hd__mux2_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07474_ _10515_/Q _07477_/S _07038_/S _07211_/X vssd1 vssd1 vccd1 vccd1 _10515_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ _11455_/Q _09206_/Y _09208_/Y _07232_/X vssd1 vssd1 vccd1 vccd1 _11455_/D
+ sky130_fd_sc_hd__o22a_1
X_06425_ _10306_/Q _08647_/B _06421_/X _06424_/X vssd1 vssd1 vccd1 vccd1 _06431_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09144_ _10171_/A1 _09132_/X _09143_/X _10175_/C1 vssd1 vssd1 vccd1 vccd1 _11417_/D
+ sky130_fd_sc_hd__o211a_1
X_06356_ _11388_/Q _09060_/A _08668_/A _11431_/Q _06355_/X vssd1 vssd1 vccd1 vccd1
+ _06356_/X sky130_fd_sc_hd__o221a_1
XFILLER_124_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05307_ _05307_/A _05307_/B _05307_/C _05307_/D vssd1 vssd1 vccd1 vccd1 _05313_/A
+ sky130_fd_sc_hd__or4_4
X_09075_ _10175_/A1 _09077_/B _08771_/A vssd1 vssd1 vccd1 vccd1 _09075_/X sky130_fd_sc_hd__a21o_1
X_06287_ _06284_/X _06286_/X _07690_/A _06282_/X vssd1 vssd1 vccd1 vccd1 _06287_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08026_ _10175_/A1 _08035_/S _08025_/X _07011_/B vssd1 vssd1 vccd1 vccd1 _10837_/D
+ sky130_fd_sc_hd__o211a_1
X_05238_ _05233_/X _05238_/B _05238_/C _05238_/D vssd1 vssd1 vccd1 vccd1 _05238_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05169_ _11224_/Q _11223_/Q _05393_/S vssd1 vssd1 vccd1 vccd1 _05176_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09977_ _09977_/A _10137_/B _10159_/C vssd1 vssd1 vccd1 vccd1 _09977_/X sky130_fd_sc_hd__or3_4
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08928_ _11323_/Q _08946_/B vssd1 vssd1 vccd1 vccd1 _08928_/X sky130_fd_sc_hd__or2_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08859_ _09275_/A1 _08884_/S _08858_/X _09092_/C1 vssd1 vssd1 vccd1 vccd1 _11286_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _11870_/A vssd1 vssd1 vccd1 vccd1 _11870_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_58_wb_clk_i clkbuf_leaf_88_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11284_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _11584_/CLK _10821_/D vssd1 vssd1 vccd1 vccd1 _10821_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10752_ _11473_/CLK _10752_/D vssd1 vssd1 vccd1 vccd1 _10752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10683_ _11703_/CLK _10683_/D vssd1 vssd1 vccd1 vccd1 _10683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11304_ _11332_/CLK _11304_/D vssd1 vssd1 vccd1 vccd1 _11304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11235_ _11235_/CLK _11235_/D vssd1 vssd1 vccd1 vccd1 _11235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11166_ _11329_/CLK _11166_/D vssd1 vssd1 vccd1 vccd1 _11166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10117_ _10117_/A0 _11764_/Q _10118_/S vssd1 vssd1 vccd1 vccd1 _11764_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11097_ _11186_/CLK _11097_/D vssd1 vssd1 vccd1 vccd1 _11097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10048_ _10058_/A _10048_/B vssd1 vssd1 vccd1 vccd1 _11715_/D sky130_fd_sc_hd__or2_1
XFILLER_75_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06210_ _06664_/C1 _06208_/X _06209_/X _06622_/A2 _05716_/X vssd1 vssd1 vccd1 vccd1
+ _06210_/X sky130_fd_sc_hd__a32o_1
X_07190_ _07190_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _07190_/X sky130_fd_sc_hd__or2_1
XFILLER_117_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06141_ _10951_/Q _06589_/A2 _06137_/X _06140_/X vssd1 vssd1 vccd1 vccd1 _06141_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06072_ _10939_/Q _06630_/A2 _06630_/B1 _11015_/Q vssd1 vssd1 vccd1 vccd1 _06072_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _11698_/Q _09566_/B _09567_/B _11713_/Q vssd1 vssd1 vccd1 vccd1 _09900_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout506 _09279_/C1 vssd1 vssd1 vccd1 vccd1 _09092_/C1 sky130_fd_sc_hd__buf_4
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout517 _08816_/A vssd1 vssd1 vccd1 vccd1 _08050_/A sky130_fd_sc_hd__buf_6
X_09831_ _09539_/B _09830_/B _09830_/Y _11587_/Q vssd1 vssd1 vccd1 vccd1 _09831_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout528 _08590_/A vssd1 vssd1 vccd1 vccd1 _08833_/A sky130_fd_sc_hd__buf_4
XFILLER_112_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout539 fanout555/X vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__buf_4
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _09515_/B _09722_/Y _09758_/Y _06955_/X vssd1 vssd1 vccd1 vccd1 _09762_/X
+ sky130_fd_sc_hd__a22o_1
X_06974_ _10221_/Q _06973_/X _09416_/A vssd1 vssd1 vccd1 vccd1 _10221_/D sky130_fd_sc_hd__mux2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08713_ _08819_/A _08713_/B vssd1 vssd1 vccd1 vccd1 _11211_/D sky130_fd_sc_hd__or2_1
X_05925_ _10875_/Q _06513_/A2 _06152_/B _10612_/Q _07083_/B vssd1 vssd1 vccd1 vccd1
+ _05925_/X sky130_fd_sc_hd__o221a_1
X_09693_ _05391_/S _09682_/B _09682_/Y _11638_/Q _09692_/X vssd1 vssd1 vccd1 vccd1
+ _09694_/B sky130_fd_sc_hd__o221a_1
XFILLER_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08644_ _11178_/Q _08645_/S _07086_/Y _08811_/B2 vssd1 vssd1 vccd1 vccd1 _11178_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05856_ _11314_/Q _09271_/A _06718_/B1 _11286_/Q _06718_/C1 vssd1 vssd1 vccd1 vccd1
+ _05856_/X sky130_fd_sc_hd__o221a_1
XFILLER_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _11143_/Q _08838_/A0 _08577_/S vssd1 vssd1 vccd1 vccd1 _08576_/B sky130_fd_sc_hd__mux2_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05787_ _11871_/A _11872_/A vssd1 vssd1 vccd1 vccd1 _05787_/X sky130_fd_sc_hd__or2_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07526_ _07930_/A _07526_/B vssd1 vssd1 vccd1 vccd1 _10547_/D sky130_fd_sc_hd__or2_1
XFILLER_74_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07457_ _10505_/Q _09226_/A _07754_/B _07456_/X vssd1 vssd1 vccd1 vccd1 _10505_/D
+ sky130_fd_sc_hd__o31a_1
X_06408_ _06535_/A _06406_/X _06407_/X _06664_/C1 vssd1 vssd1 vccd1 vccd1 _06408_/X
+ sky130_fd_sc_hd__o211a_1
X_07388_ _10470_/Q _10132_/A0 _07393_/S vssd1 vssd1 vccd1 vccd1 _07389_/B sky130_fd_sc_hd__mux2_1
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09127_ _11410_/Q _09127_/B vssd1 vssd1 vccd1 vccd1 _09127_/X sky130_fd_sc_hd__or2_1
X_06339_ _07689_/A _06337_/X _06338_/X _07082_/A vssd1 vssd1 vccd1 vccd1 _06339_/X
+ sky130_fd_sc_hd__a211o_4
Xclkbuf_leaf_105_wb_clk_i clkbuf_4_10__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11450_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09058_ _11378_/Q _09038_/X _09057_/X vssd1 vssd1 vccd1 vccd1 _11378_/D sky130_fd_sc_hd__a21o_1
XFILLER_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08009_ _07061_/A _10829_/Q _08011_/S vssd1 vssd1 vccd1 vccd1 _08010_/B sky130_fd_sc_hd__mux2_1
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11020_ _11312_/CLK _11020_/D vssd1 vssd1 vccd1 vccd1 _11020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1120 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1120/HI irq[0] sky130_fd_sc_hd__conb_1
XFILLER_46_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1131 vssd1 vssd1 vccd1 vccd1 io_oeb[8] wrapped_tms1x00_1131/LO sky130_fd_sc_hd__conb_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10804_ _10804_/CLK _10804_/D vssd1 vssd1 vccd1 vccd1 _10804_/Q sky130_fd_sc_hd__dfxtp_1
X_11784_ _11791_/CLK _11784_/D vssd1 vssd1 vccd1 vccd1 _11784_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10735_ _10735_/CLK _10735_/D vssd1 vssd1 vccd1 vccd1 _10735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10666_ _10666_/CLK _10666_/D vssd1 vssd1 vccd1 vccd1 _10666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10597_ _11768_/CLK _10597_/D vssd1 vssd1 vccd1 vccd1 _10597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11218_ _11220_/CLK _11218_/D vssd1 vssd1 vccd1 vccd1 _11218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11149_ _11151_/CLK _11149_/D vssd1 vssd1 vccd1 vccd1 _11149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05710_ _11038_/Q _05609_/Y _05627_/Y _11033_/Q vssd1 vssd1 vccd1 vccd1 _05710_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06690_ _10710_/Q _07778_/A _06727_/B _10408_/Q vssd1 vssd1 vccd1 vccd1 _06690_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_64_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05641_ _11329_/Q _05579_/Y _05597_/Y _11320_/Q vssd1 vssd1 vccd1 vccd1 _05641_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08360_ _08838_/A0 _11023_/Q _08360_/S vssd1 vssd1 vccd1 vccd1 _08361_/B sky130_fd_sc_hd__mux2_1
X_05572_ _05076_/A _11418_/Q _11413_/Q _05620_/B2 _05571_/X vssd1 vssd1 vccd1 vccd1
+ _05573_/B sky130_fd_sc_hd__a221o_4
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11777_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07311_ _10421_/Q _07301_/Y _07306_/Y _07016_/X vssd1 vssd1 vccd1 vccd1 _10421_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08291_ _10977_/Q _07090_/X _08298_/S vssd1 vssd1 vccd1 vccd1 _10977_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07242_ _07241_/X _10389_/Q _07249_/S vssd1 vssd1 vccd1 vccd1 _10389_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07173_ _07920_/A _07173_/B vssd1 vssd1 vccd1 vccd1 _10347_/D sky130_fd_sc_hd__or2_1
XFILLER_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06124_ _10460_/Q _06308_/A2 _10009_/A _11308_/Q _06123_/X vssd1 vssd1 vccd1 vccd1
+ _06125_/C sky130_fd_sc_hd__o221a_1
XFILLER_118_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06055_ _11127_/Q _06635_/A2 _06556_/B1 _10302_/Q vssd1 vssd1 vccd1 vccd1 _06055_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout303 _07557_/S vssd1 vssd1 vccd1 vccd1 _07593_/S sky130_fd_sc_hd__buf_6
Xfanout314 _07440_/X vssd1 vssd1 vccd1 vccd1 _07535_/S sky130_fd_sc_hd__buf_8
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout325 _07202_/Y vssd1 vssd1 vccd1 vccd1 _07204_/B sky130_fd_sc_hd__buf_12
XFILLER_87_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout336 _07045_/Y vssd1 vssd1 vccd1 vccd1 _07078_/B sky130_fd_sc_hd__buf_6
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09814_ _10529_/Q _09572_/B _09566_/D _10531_/Q _09801_/X vssd1 vssd1 vccd1 vccd1
+ _09815_/D sky130_fd_sc_hd__a221o_1
Xfanout347 _07102_/X vssd1 vssd1 vccd1 vccd1 _08901_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout358 _10159_/B vssd1 vssd1 vccd1 vccd1 _09271_/B sky130_fd_sc_hd__buf_8
XFILLER_28_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout369 _08323_/A vssd1 vssd1 vccd1 vccd1 _08437_/A sky130_fd_sc_hd__buf_6
XFILLER_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09745_ _10537_/Q _09877_/A2 _09875_/A2 _10497_/Q vssd1 vssd1 vccd1 vccd1 _09745_/X
+ sky130_fd_sc_hd__a22o_1
X_06957_ input7/X _09538_/D _06956_/Y _06950_/A vssd1 vssd1 vccd1 vccd1 _06957_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05908_ _10620_/Q _07222_/A _06105_/B1 _10718_/Q vssd1 vssd1 vccd1 vccd1 _05908_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ _07007_/A _07048_/A _08970_/S _06884_/Y _10214_/Q vssd1 vssd1 vccd1 vccd1
+ _10214_/D sky130_fd_sc_hd__a32o_1
X_09676_ _09672_/Y _09674_/Y _09554_/Y vssd1 vssd1 vccd1 vccd1 _09676_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05839_ _10257_/Q _06976_/A _06903_/A _10194_/Q vssd1 vssd1 vccd1 vccd1 _05839_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08627_ _11168_/Q _08633_/B vssd1 vssd1 vccd1 vccd1 _08627_/X sky130_fd_sc_hd__or2_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08558_ _11134_/Q _10135_/A0 _08558_/S vssd1 vssd1 vccd1 vccd1 _08559_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07509_ _08929_/A1 _10539_/Q _07533_/S vssd1 vssd1 vccd1 vccd1 _07510_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08489_ _11095_/Q _08503_/B vssd1 vssd1 vccd1 vccd1 _08489_/X sky130_fd_sc_hd__or2_1
XFILLER_74_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10520_ _11711_/CLK _10520_/D vssd1 vssd1 vccd1 vccd1 _10520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10451_ _11310_/CLK _10451_/D vssd1 vssd1 vccd1 vccd1 _10451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10382_ _11702_/CLK _10382_/D vssd1 vssd1 vccd1 vccd1 _10382_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_100_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11003_ _11005_/CLK _11003_/D vssd1 vssd1 vccd1 vccd1 _11003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_73_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11495_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout870 _06719_/A2 vssd1 vssd1 vccd1 vccd1 _06455_/A2 sky130_fd_sc_hd__buf_6
XFILLER_120_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout881 _06553_/B vssd1 vssd1 vccd1 vccd1 _06370_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout892 _06194_/A2 vssd1 vssd1 vccd1 vccd1 _06862_/A2 sky130_fd_sc_hd__buf_8
XFILLER_93_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11777_/CLK _11767_/D vssd1 vssd1 vccd1 vccd1 _11767_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10718_ _10727_/CLK _10718_/D vssd1 vssd1 vccd1 vccd1 _10718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11698_ _11698_/CLK _11698_/D vssd1 vssd1 vccd1 vccd1 _11698_/Q sky130_fd_sc_hd__dfxtp_1
X_10649_ _11270_/CLK _10649_/D vssd1 vssd1 vccd1 vccd1 _10649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07860_ _10015_/A0 _07871_/S _07859_/X _07868_/C1 vssd1 vssd1 vccd1 vccd1 _10748_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06811_ _06577_/A _10246_/Q _06853_/A3 _06810_/X _05730_/Y vssd1 vssd1 vccd1 vccd1
+ _06811_/X sky130_fd_sc_hd__a32o_1
X_07791_ _10021_/A0 _10703_/Q _09193_/B vssd1 vssd1 vccd1 vccd1 _07792_/B sky130_fd_sc_hd__mux2_1
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06742_ _11619_/Q _06741_/X _06883_/B vssd1 vssd1 vccd1 vccd1 _10241_/D sky130_fd_sc_hd__mux2_1
X_09530_ _09492_/B _09522_/B _09504_/B _09489_/C _11620_/Q vssd1 vssd1 vccd1 vccd1
+ _09530_/X sky130_fd_sc_hd__a41o_1
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09461_ input36/X _09442_/X _09460_/X vssd1 vssd1 vccd1 vccd1 _09462_/B sky130_fd_sc_hd__o21ai_1
X_06673_ _10758_/Q _07854_/A _06806_/A2 _10570_/Q _06672_/X vssd1 vssd1 vccd1 vccd1
+ _06673_/X sky130_fd_sc_hd__o221a_1
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05624_ _11749_/Q _05630_/A2 _05630_/B1 _11747_/Q _05622_/X vssd1 vssd1 vccd1 vccd1
+ _05627_/A sky130_fd_sc_hd__a221o_4
XFILLER_58_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08412_ _09182_/A0 _11047_/Q _08414_/S vssd1 vssd1 vccd1 vccd1 _08413_/B sky130_fd_sc_hd__mux2_1
X_09392_ _09999_/A0 _11558_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _11558_/D sky130_fd_sc_hd__mux2_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08343_ _08492_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _11014_/D sky130_fd_sc_hd__or2_1
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05555_ _05555_/A _05555_/B vssd1 vssd1 vccd1 vccd1 _05555_/Y sky130_fd_sc_hd__nor2_8
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08274_ _09182_/A0 _10969_/Q _08276_/S vssd1 vssd1 vccd1 vccd1 _08275_/B sky130_fd_sc_hd__mux2_1
X_05486_ _10231_/Q input73/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05486_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07225_ _07225_/A _08322_/A vssd1 vssd1 vccd1 vccd1 _07225_/X sky130_fd_sc_hd__or2_4
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07156_ _10013_/A0 _10339_/Q _09243_/C vssd1 vssd1 vccd1 vccd1 _07157_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06107_ _10686_/Q _07904_/A _06857_/B1 _11700_/Q vssd1 vssd1 vccd1 vccd1 _06107_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07087_ _08819_/A _08645_/S vssd1 vssd1 vccd1 vccd1 _07109_/S sky130_fd_sc_hd__or2_4
XFILLER_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06038_ _10207_/Q _06351_/A2 _06034_/X _06037_/X vssd1 vssd1 vccd1 vccd1 _06038_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07989_ _10820_/Q _08818_/A1 _07991_/S vssd1 vssd1 vccd1 vccd1 _07990_/B sky130_fd_sc_hd__mux2_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09728_ _10346_/Q _09884_/A2 _09565_/C _11468_/Q _09727_/X vssd1 vssd1 vccd1 vccd1
+ _09731_/C sky130_fd_sc_hd__a221o_1
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09659_ _09659_/A _09659_/B _09659_/C _09659_/D vssd1 vssd1 vccd1 vccd1 _09659_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11621_ _11812_/CLK _11621_/D vssd1 vssd1 vccd1 vccd1 _11621_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_120_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11745_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11552_ _11675_/CLK _11552_/D vssd1 vssd1 vccd1 vccd1 _11552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10503_ _11450_/CLK _10503_/D vssd1 vssd1 vccd1 vccd1 _10503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11483_ _11809_/CLK _11483_/D vssd1 vssd1 vccd1 vccd1 _11483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10434_ _11284_/CLK _10434_/D vssd1 vssd1 vccd1 vccd1 _10434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10365_ _10798_/CLK _10365_/D vssd1 vssd1 vccd1 vccd1 _10365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _11716_/CLK _10296_/D vssd1 vssd1 vccd1 vccd1 _10296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05340_ _05340_/A _05340_/B _05340_/C _05340_/D vssd1 vssd1 vccd1 vccd1 _05346_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05271_ _10454_/Q _10453_/Q _05385_/S vssd1 vssd1 vccd1 vccd1 _05275_/A sky130_fd_sc_hd__mux2_1
X_07010_ _07010_/A _10028_/A vssd1 vssd1 vccd1 vccd1 _07227_/B sky130_fd_sc_hd__and2_4
XFILLER_122_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08961_ _08965_/A _08961_/B vssd1 vssd1 vccd1 vccd1 _08961_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07912_ _07926_/A _07912_/B vssd1 vssd1 vccd1 vccd1 _10773_/D sky130_fd_sc_hd__or2_1
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08892_ _11303_/Q _08894_/B vssd1 vssd1 vccd1 vccd1 _08892_/X sky130_fd_sc_hd__or2_1
XFILLER_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07843_ _09232_/B2 _10738_/Q _07846_/S vssd1 vssd1 vccd1 vccd1 _10738_/D sky130_fd_sc_hd__mux2_1
XFILLER_151_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07774_ _10051_/A1 _07776_/A2 _07204_/Y _10694_/Q _07451_/A vssd1 vssd1 vccd1 vccd1
+ _10694_/D sky130_fd_sc_hd__a221o_1
X_09513_ _09525_/A _09500_/B _09512_/A _11614_/Q vssd1 vssd1 vccd1 vccd1 _09513_/X
+ sky130_fd_sc_hd__a31o_1
X_06725_ _11714_/Q _10009_/A _07819_/A _10800_/Q _06724_/X vssd1 vssd1 vccd1 vccd1
+ _06725_/X sky130_fd_sc_hd__o221a_1
XFILLER_65_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09444_ _09444_/A _09478_/A vssd1 vssd1 vccd1 vccd1 _09444_/Y sky130_fd_sc_hd__nand2_1
X_06656_ _11048_/Q _05736_/Y _05746_/X _10970_/Q vssd1 vssd1 vccd1 vccd1 _06656_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05607_ _05631_/A2 _11547_/Q _11543_/Q _05631_/B1 _05605_/X vssd1 vssd1 vccd1 vccd1
+ _05607_/X sky130_fd_sc_hd__a221o_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ _10175_/A1 _09359_/X _09374_/X _09995_/C1 vssd1 vssd1 vccd1 vccd1 _11545_/D
+ sky130_fd_sc_hd__o211a_1
X_06587_ _11277_/Q _06628_/B1 _06630_/B1 _11023_/Q vssd1 vssd1 vccd1 vccd1 _06587_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05538_ _05628_/A2 _11356_/Q _11353_/Q _05628_/B1 vssd1 vssd1 vccd1 vccd1 _05538_/X
+ sky130_fd_sc_hd__a22o_1
X_08326_ _11001_/Q _08322_/Y _08325_/Y _08326_/B2 vssd1 vssd1 vccd1 vccd1 _11001_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_138_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08257_ _08869_/A _08257_/B vssd1 vssd1 vccd1 vccd1 _10960_/D sky130_fd_sc_hd__or2_1
X_05469_ _05469_/A _05469_/B _05469_/C _05469_/D vssd1 vssd1 vccd1 vccd1 _05470_/B
+ sky130_fd_sc_hd__or4_1
X_07208_ _07057_/A _07204_/B _07771_/B1 _10366_/Q vssd1 vssd1 vccd1 vccd1 _10366_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08188_ _10928_/Q _08197_/S _07644_/Y _08811_/B2 vssd1 vssd1 vccd1 vccd1 _10928_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07139_ _10331_/Q _07145_/B vssd1 vssd1 vccd1 vccd1 _07139_/X sky130_fd_sc_hd__or2_1
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10150_ _10150_/A1 _10154_/B _10150_/B1 vssd1 vssd1 vccd1 vccd1 _10150_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10081_ _10117_/A0 _11741_/Q _10082_/S vssd1 vssd1 vccd1 vccd1 _11741_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10983_ _11310_/CLK _10983_/D vssd1 vssd1 vccd1 vccd1 _10983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11604_ _11604_/CLK _11604_/D vssd1 vssd1 vccd1 vccd1 _11604_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_141_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11535_ _11735_/CLK _11535_/D vssd1 vssd1 vccd1 vccd1 _11535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11466_ _11471_/CLK _11466_/D vssd1 vssd1 vccd1 vccd1 _11466_/Q sky130_fd_sc_hd__dfxtp_2
X_10417_ _10644_/CLK _10417_/D vssd1 vssd1 vccd1 vccd1 _10417_/Q sky130_fd_sc_hd__dfxtp_1
X_11397_ _11410_/CLK _11397_/D vssd1 vssd1 vccd1 vccd1 _11397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10348_ _11462_/CLK _10348_/D vssd1 vssd1 vccd1 vccd1 _10348_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10279_ _11745_/CLK _10279_/D vssd1 vssd1 vccd1 vccd1 _10279_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06510_ _10818_/Q _06639_/B1 _06506_/X _06509_/X vssd1 vssd1 vccd1 vccd1 _06510_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07490_ _07108_/X _10526_/Q _07490_/S vssd1 vssd1 vccd1 vccd1 _10526_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06441_ _11705_/Q _08560_/A _06438_/X _06440_/X vssd1 vssd1 vccd1 vccd1 _06441_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_22_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09160_ _09364_/A1 _09154_/X _09159_/X _10175_/C1 vssd1 vssd1 vccd1 vccd1 _11424_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06372_ _10483_/Q _07190_/A _10009_/A _11704_/Q _06550_/C1 vssd1 vssd1 vccd1 vccd1
+ _06374_/B sky130_fd_sc_hd__o221a_1
X_08111_ _10881_/Q _10128_/A0 _08120_/S vssd1 vssd1 vccd1 vccd1 _08112_/B sky130_fd_sc_hd__mux2_1
X_05323_ _05323_/A _05323_/B _05323_/C _05323_/D vssd1 vssd1 vccd1 vccd1 _05324_/B
+ sky130_fd_sc_hd__or4_4
X_09091_ _11393_/Q _09099_/B vssd1 vssd1 vccd1 vccd1 _09091_/X sky130_fd_sc_hd__or2_1
XFILLER_30_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08042_ _10846_/Q _10128_/A0 _08051_/S vssd1 vssd1 vccd1 vccd1 _08043_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05254_ _10984_/Q _10983_/Q _05385_/S vssd1 vssd1 vccd1 vccd1 _05258_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05185_ _10834_/Q _10591_/Q _09539_/B vssd1 vssd1 vccd1 vccd1 _05189_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ _10175_/A1 _09977_/X _09992_/X _09993_/C1 vssd1 vssd1 vccd1 vccd1 _11683_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ _11331_/Q _08946_/B vssd1 vssd1 vccd1 vccd1 _08944_/X sky130_fd_sc_hd__or2_1
XFILLER_130_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08875_ _08875_/A _08875_/B vssd1 vssd1 vccd1 vccd1 _11294_/D sky130_fd_sc_hd__or2_1
XFILLER_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07826_ _09214_/A _07820_/B _07956_/S _10721_/Q vssd1 vssd1 vccd1 vccd1 _10721_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07757_ _07036_/A _07761_/A2 _07756_/X _09201_/A1 vssd1 vssd1 vccd1 vccd1 _10679_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06708_ _10409_/Q _06727_/B _06707_/X _06878_/C1 vssd1 vssd1 vccd1 vccd1 _06708_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07688_ _10644_/Q _07674_/X _07675_/Y _07318_/X vssd1 vssd1 vccd1 vccd1 _10644_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_73_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ _11634_/Q _11586_/Q _09704_/B vssd1 vssd1 vccd1 vccd1 _11586_/D sky130_fd_sc_hd__mux2_1
X_06639_ _10887_/Q _06553_/B _06639_/B1 _10821_/Q vssd1 vssd1 vccd1 vccd1 _06639_/X
+ sky130_fd_sc_hd__o22a_1
X_09358_ _09358_/A _10158_/B _10158_/C vssd1 vssd1 vccd1 vccd1 _09376_/B sky130_fd_sc_hd__and3_4
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08309_ _10989_/Q _08302_/Y _08303_/Y _07095_/X vssd1 vssd1 vccd1 vccd1 _10989_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_138_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09289_ _09289_/A1 _09271_/X _09288_/X _09289_/C1 vssd1 vssd1 vccd1 vccd1 _11496_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11320_ _11330_/CLK _11320_/D vssd1 vssd1 vccd1 vccd1 _11320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11251_ _11251_/CLK _11251_/D vssd1 vssd1 vccd1 vccd1 _11251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10202_ _11803_/CLK _10202_/D vssd1 vssd1 vccd1 vccd1 _10202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ _11224_/CLK _11182_/D vssd1 vssd1 vccd1 vccd1 _11182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10133_ _08661_/A _11779_/Q _10135_/S vssd1 vssd1 vccd1 vccd1 _11779_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10064_ _10111_/A0 _11725_/Q _10071_/S vssd1 vssd1 vccd1 vccd1 _11725_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10966_ _11683_/CLK _10966_/D vssd1 vssd1 vccd1 vccd1 _10966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10897_ _11601_/CLK _10897_/D vssd1 vssd1 vccd1 vccd1 _10897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11518_ _11683_/CLK _11518_/D vssd1 vssd1 vccd1 vccd1 _11518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11449_ _11462_/CLK _11449_/D vssd1 vssd1 vccd1 vccd1 _11449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06990_ _10150_/A1 _06976_/X _06989_/X _06990_/C1 vssd1 vssd1 vccd1 vccd1 _10262_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05941_ _11055_/Q _06631_/A2 _08123_/A _10889_/Q _06392_/C1 vssd1 vssd1 vccd1 vccd1
+ _05941_/X sky130_fd_sc_hd__o221a_1
XFILLER_152_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05872_ _10787_/Q _06455_/A2 _06412_/B1 _10834_/Q vssd1 vssd1 vccd1 vccd1 _05872_/X
+ sky130_fd_sc_hd__o22a_1
X_08660_ _08757_/A _08660_/B vssd1 vssd1 vccd1 vccd1 _11185_/D sky130_fd_sc_hd__or2_1
XFILLER_27_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07611_ _09037_/A _08471_/B _10136_/C vssd1 vssd1 vccd1 vccd1 _08037_/B sky130_fd_sc_hd__and3_4
X_08591_ _11151_/Q _08591_/B vssd1 vssd1 vccd1 vccd1 _08591_/X sky130_fd_sc_hd__or2_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07542_ _08781_/A _07542_/B vssd1 vssd1 vccd1 vccd1 _10554_/D sky130_fd_sc_hd__or2_1
XFILLER_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07473_ _07476_/A _07473_/B vssd1 vssd1 vccd1 vccd1 _10514_/D sky130_fd_sc_hd__or2_1
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09212_ _11454_/Q _09206_/Y _09208_/Y _07093_/X vssd1 vssd1 vccd1 vccd1 _11454_/D
+ sky130_fd_sc_hd__o22a_1
X_06424_ _10598_/Q _06731_/B1 _06423_/X _11869_/A vssd1 vssd1 vccd1 vccd1 _06424_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09143_ _11417_/Q _09149_/B vssd1 vssd1 vccd1 vccd1 _09143_/X sky130_fd_sc_hd__or2_1
X_06355_ _11497_/Q _09271_/A _08972_/A _11348_/Q vssd1 vssd1 vccd1 vccd1 _06355_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_33_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05306_ _11016_/Q _11015_/Q _05372_/S vssd1 vssd1 vccd1 vccd1 _05307_/D sky130_fd_sc_hd__mux2_1
X_09074_ _09285_/A1 _09060_/X _09073_/X _09078_/C1 vssd1 vssd1 vccd1 vccd1 _11385_/D
+ sky130_fd_sc_hd__o211a_1
X_06286_ _10264_/Q _06976_/A _06351_/A2 _10211_/Q _06285_/X vssd1 vssd1 vccd1 vccd1
+ _06286_/X sky130_fd_sc_hd__o221a_1
XFILLER_136_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08025_ _10837_/Q _08037_/B vssd1 vssd1 vccd1 vccd1 _08025_/X sky130_fd_sc_hd__or2_1
X_05237_ _05237_/A _05237_/B vssd1 vssd1 vccd1 vccd1 _05238_/D sky130_fd_sc_hd__nor2_1
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05168_ _05168_/A _05168_/B vssd1 vssd1 vccd1 vccd1 _05168_/Y sky130_fd_sc_hd__nor2_2
XFILLER_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09976_ _09976_/A _10158_/B _10158_/C vssd1 vssd1 vccd1 vccd1 _09994_/B sky130_fd_sc_hd__and3_4
X_05099_ _11577_/Q vssd1 vssd1 vccd1 vccd1 _09441_/B sky130_fd_sc_hd__inv_2
XFILLER_103_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08927_ _09101_/A1 _08945_/A2 _08926_/X _08947_/C1 vssd1 vssd1 vccd1 vccd1 _11322_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08858_ _11286_/Q _08894_/B vssd1 vssd1 vccd1 vccd1 _08858_/X sky130_fd_sc_hd__or2_1
XFILLER_40_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07809_ _07932_/A1 _10712_/Q _09193_/B vssd1 vssd1 vccd1 vccd1 _07810_/B sky130_fd_sc_hd__mux2_1
XFILLER_57_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ _08789_/A1 _08792_/S _08788_/X _09168_/C1 vssd1 vssd1 vccd1 vccd1 _11250_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _11584_/CLK _10820_/D vssd1 vssd1 vccd1 vccd1 _10820_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_98_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _10666_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10751_ _11622_/CLK _10751_/D vssd1 vssd1 vccd1 vccd1 _10751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11604_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10682_ _11698_/CLK _10682_/D vssd1 vssd1 vccd1 vccd1 _10682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11303_ _11393_/CLK _11303_/D vssd1 vssd1 vccd1 vccd1 _11303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11234_ _11234_/CLK _11234_/D vssd1 vssd1 vccd1 vccd1 _11234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11165_ _11243_/CLK _11165_/D vssd1 vssd1 vccd1 vccd1 _11165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10116_ _07018_/A _11763_/Q _10118_/S vssd1 vssd1 vccd1 vccd1 _11763_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11096_ _11312_/CLK _11096_/D vssd1 vssd1 vccd1 vccd1 _11096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10047_ _11715_/Q _10047_/A1 _10057_/S vssd1 vssd1 vccd1 vccd1 _10048_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10949_ _11235_/CLK _10949_/D vssd1 vssd1 vccd1 vccd1 _10949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06140_ _11280_/Q _06227_/A2 _06139_/X _06265_/C1 vssd1 vssd1 vccd1 vccd1 _06140_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06071_ _11057_/Q _08054_/A _08123_/A _10891_/Q _06392_/C1 vssd1 vssd1 vccd1 vccd1
+ _06071_/X sky130_fd_sc_hd__o221a_1
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09830_ _11657_/Q _09830_/B vssd1 vssd1 vccd1 vccd1 _09830_/Y sky130_fd_sc_hd__nand2_1
Xfanout507 _09279_/C1 vssd1 vssd1 vccd1 vccd1 _08919_/C1 sky130_fd_sc_hd__clkbuf_4
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout518 _07659_/A vssd1 vssd1 vccd1 vccd1 _08816_/A sky130_fd_sc_hd__buf_4
XFILLER_99_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout529 _08492_/A vssd1 vssd1 vccd1 vccd1 _08590_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _11643_/Q _09760_/X _09770_/S vssd1 vssd1 vccd1 vccd1 _11643_/D sky130_fd_sc_hd__mux2_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _11665_/Q _05474_/B _06969_/X _05474_/A _06972_/X vssd1 vssd1 vccd1 vccd1
+ _06973_/X sky130_fd_sc_hd__a221o_4
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _11211_/Q _07092_/A _08726_/S vssd1 vssd1 vccd1 vccd1 _08713_/B sky130_fd_sc_hd__mux2_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05924_ _10457_/Q _06308_/A2 _07111_/A _10810_/Q vssd1 vssd1 vccd1 vccd1 _05924_/X
+ sky130_fd_sc_hd__o22a_1
X_09692_ _11642_/Q _09692_/B vssd1 vssd1 vccd1 vccd1 _09692_/X sky130_fd_sc_hd__or2_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08643_ _11177_/Q _08645_/S _07086_/Y _07617_/B vssd1 vssd1 vccd1 vccd1 _11177_/D
+ sky130_fd_sc_hd__o22a_1
X_05855_ _11190_/Q _06719_/A2 _06716_/B1 _11240_/Q vssd1 vssd1 vccd1 vccd1 _05855_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ _11142_/Q _08577_/S _08563_/Y _08817_/B2 vssd1 vssd1 vccd1 vccd1 _11142_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05786_ _11871_/A _11872_/A vssd1 vssd1 vccd1 vccd1 _05786_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ _07932_/A1 _10547_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _07526_/B sky130_fd_sc_hd__mux2_1
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07456_ _10015_/A0 _07441_/A _07755_/A2 _09241_/B1 vssd1 vssd1 vccd1 vccd1 _07456_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06407_ _06382_/X _06405_/X _06576_/A vssd1 vssd1 vccd1 vccd1 _06407_/X sky130_fd_sc_hd__a21o_1
X_07387_ _10469_/Q _07393_/S _07655_/S _07098_/B vssd1 vssd1 vccd1 vccd1 _10469_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09126_ _11409_/Q _09110_/X _09125_/X vssd1 vssd1 vccd1 vccd1 _11409_/D sky130_fd_sc_hd__a21o_1
XFILLER_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06338_ _06322_/X _06327_/X _07690_/A vssd1 vssd1 vccd1 vccd1 _06338_/X sky130_fd_sc_hd__o21a_1
XFILLER_136_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09057_ _10178_/A1 _09055_/B _09173_/B1 vssd1 vssd1 vccd1 vccd1 _09057_/X sky130_fd_sc_hd__a21o_1
X_06269_ _11312_/Q _06459_/A2 _06459_/B1 _10874_/Q vssd1 vssd1 vccd1 vccd1 _06269_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ _07059_/A _08015_/S _08007_/X _08831_/C1 vssd1 vssd1 vccd1 vccd1 _10828_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09959_ _09959_/A _09959_/B _09959_/C vssd1 vssd1 vccd1 vccd1 _09963_/B sky130_fd_sc_hd__nor3_4
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_tms1x00_1110 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1110/HI io_out[2] sky130_fd_sc_hd__conb_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1121 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1121/HI irq[1] sky130_fd_sc_hd__conb_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1132 vssd1 vssd1 vccd1 vccd1 io_oeb[9] wrapped_tms1x00_1132/LO sky130_fd_sc_hd__conb_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10803_ _11474_/CLK _10803_/D vssd1 vssd1 vccd1 vccd1 _10803_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _11809_/CLK _11783_/D vssd1 vssd1 vccd1 vccd1 _11783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10734_ _11722_/CLK _10734_/D vssd1 vssd1 vccd1 vccd1 _10734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10665_ _11457_/CLK _10665_/D vssd1 vssd1 vccd1 vccd1 _10665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10596_ _11284_/CLK _10596_/D vssd1 vssd1 vccd1 vccd1 _10596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11217_ _11220_/CLK _11217_/D vssd1 vssd1 vccd1 vccd1 _11217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11148_ _11151_/CLK _11148_/D vssd1 vssd1 vccd1 vccd1 _11148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11079_ _11781_/CLK _11079_/D vssd1 vssd1 vccd1 vccd1 _11079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05640_ _11321_/Q _05549_/Y _05555_/Y _11324_/Q _05639_/X vssd1 vssd1 vccd1 vccd1
+ _05643_/B sky130_fd_sc_hd__a221o_1
XFILLER_24_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05571_ _05619_/A1 _11421_/Q _11417_/Q _05619_/B2 _05568_/X vssd1 vssd1 vccd1 vccd1
+ _05571_/X sky130_fd_sc_hd__a221o_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07310_ _10420_/Q _07302_/Y _07305_/Y _07309_/X vssd1 vssd1 vccd1 vccd1 _10420_/D
+ sky130_fd_sc_hd__o22a_1
X_08290_ _10976_/Q _08326_/B2 _08298_/S vssd1 vssd1 vccd1 vccd1 _10976_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07241_ _07451_/A _07241_/B vssd1 vssd1 vccd1 vccd1 _07241_/X sky130_fd_sc_hd__or2_1
XFILLER_121_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07172_ _08883_/A1 _10347_/Q _07172_/S vssd1 vssd1 vccd1 vccd1 _07173_/B sky130_fd_sc_hd__mux2_1
XFILLER_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06123_ _10465_/Q _06371_/A2 _07827_/A2 _10980_/Q vssd1 vssd1 vccd1 vccd1 _06123_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_8_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06054_ _11107_/Q _06539_/A2 _06050_/X _06053_/X vssd1 vssd1 vccd1 vccd1 _06054_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_105_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout304 _07557_/S vssd1 vssd1 vccd1 vccd1 _07589_/S sky130_fd_sc_hd__buf_6
XFILLER_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout315 _07380_/S vssd1 vssd1 vccd1 vccd1 _07393_/S sky130_fd_sc_hd__buf_12
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout326 _07202_/Y vssd1 vssd1 vccd1 vccd1 _07776_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout337 _07045_/Y vssd1 vssd1 vccd1 vccd1 _07047_/B sky130_fd_sc_hd__buf_6
X_09813_ _10293_/Q _09567_/B _09944_/B1 _10291_/Q _09806_/X vssd1 vssd1 vccd1 vccd1
+ _09815_/C sky130_fd_sc_hd__a221o_1
XFILLER_99_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout348 _08665_/C vssd1 vssd1 vccd1 vccd1 _10119_/B sky130_fd_sc_hd__buf_6
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout359 _10136_/B vssd1 vssd1 vccd1 vccd1 _10158_/B sky130_fd_sc_hd__buf_6
XFILLER_45_1370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09744_ _10534_/Q _09873_/A2 _09567_/C _10538_/Q _09743_/X vssd1 vssd1 vccd1 vccd1
+ _09749_/B sky130_fd_sc_hd__a221o_1
XFILLER_74_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06956_ _08956_/B _09538_/D vssd1 vssd1 vccd1 vccd1 _06956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05907_ _05891_/X _05896_/X _05906_/X _06189_/A1 vssd1 vssd1 vccd1 vccd1 _05907_/X
+ sky130_fd_sc_hd__o22a_1
X_09675_ _11633_/Q _09672_/Y _09674_/Y _11632_/Q vssd1 vssd1 vccd1 vccd1 _09675_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06887_ _07002_/A _07048_/A _08970_/S _06884_/Y _10215_/Q vssd1 vssd1 vccd1 vccd1
+ _10215_/D sky130_fd_sc_hd__a32o_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08626_ _08853_/A1 _08623_/S _08625_/X _08937_/C1 vssd1 vssd1 vccd1 vccd1 _11167_/D
+ sky130_fd_sc_hd__o211a_1
X_05838_ _11360_/Q _09016_/A _08994_/A _11350_/Q _06349_/C1 vssd1 vssd1 vccd1 vccd1
+ _05838_/X sky130_fd_sc_hd__o221a_1
XFILLER_82_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _11133_/Q _07353_/B _07357_/S _07333_/B vssd1 vssd1 vccd1 vccd1 _11133_/D
+ sky130_fd_sc_hd__o22a_1
X_05769_ _11359_/Q _10087_/A _10137_/A _11349_/Q _06214_/C1 vssd1 vssd1 vccd1 vccd1
+ _05769_/X sky130_fd_sc_hd__o221a_1
X_07508_ _09129_/A1 _07533_/S _07507_/X _07866_/C1 vssd1 vssd1 vccd1 vccd1 _10538_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08488_ _08833_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _11094_/D sky130_fd_sc_hd__or2_1
XFILLER_126_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07439_ _07440_/A _07854_/B vssd1 vssd1 vccd1 vccd1 _07537_/B sky130_fd_sc_hd__nor2_8
XFILLER_52_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10450_ _11780_/CLK _10450_/D vssd1 vssd1 vccd1 vccd1 _10450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09109_ _09109_/A _10136_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09127_/B sky130_fd_sc_hd__and3_4
XFILLER_109_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10381_ _11713_/CLK _10381_/D vssd1 vssd1 vccd1 vccd1 _10381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ _11234_/CLK _11002_/D vssd1 vssd1 vccd1 vccd1 _11002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout860 fanout861/X vssd1 vssd1 vccd1 vccd1 _06230_/A2 sky130_fd_sc_hd__buf_4
XFILLER_77_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout871 _06736_/A2 vssd1 vssd1 vccd1 vccd1 _08668_/A sky130_fd_sc_hd__buf_6
Xfanout882 _06631_/A2 vssd1 vssd1 vccd1 vccd1 _08054_/A sky130_fd_sc_hd__buf_4
Xfanout893 fanout901/X vssd1 vssd1 vccd1 vccd1 _06194_/A2 sky130_fd_sc_hd__buf_8
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11808_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11766_ _11766_/CLK _11766_/D vssd1 vssd1 vccd1 vccd1 _11766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ _10725_/CLK _10717_/D vssd1 vssd1 vccd1 vccd1 _10717_/Q sky130_fd_sc_hd__dfxtp_1
X_11697_ _11698_/CLK _11697_/D vssd1 vssd1 vccd1 vccd1 _11697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10648_ _11270_/CLK _10648_/D vssd1 vssd1 vccd1 vccd1 _10648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10579_ _11477_/CLK _10579_/D vssd1 vssd1 vccd1 vccd1 _10579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06810_ _06577_/A _10246_/Q _06852_/A3 _06743_/X _06809_/X vssd1 vssd1 vccd1 vccd1
+ _06810_/X sky130_fd_sc_hd__a32o_1
X_07790_ _07790_/A _07790_/B vssd1 vssd1 vccd1 vccd1 _10702_/D sky130_fd_sc_hd__or2_1
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06741_ _05734_/X _06734_/X _06739_/X _06740_/X vssd1 vssd1 vccd1 vccd1 _06741_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09460_ _09441_/A input22/X _09441_/Y input30/X _09459_/X vssd1 vssd1 vccd1 vccd1
+ _09460_/X sky130_fd_sc_hd__a221o_1
XFILLER_149_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06672_ _11457_/Q _06875_/A2 _06766_/A2 _11469_/Q vssd1 vssd1 vccd1 vccd1 _06672_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_64_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08411_ _08935_/A1 _08414_/S _08410_/X _07003_/B vssd1 vssd1 vccd1 vccd1 _11046_/D
+ sky130_fd_sc_hd__o211a_1
X_05623_ _11754_/Q _05629_/A2 _05629_/B1 _11748_/Q vssd1 vssd1 vccd1 vccd1 _05623_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09391_ _09391_/A _10180_/B _10180_/C vssd1 vssd1 vccd1 vccd1 _09401_/S sky130_fd_sc_hd__or3_4
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08342_ _10112_/A0 _11014_/Q _08360_/S vssd1 vssd1 vccd1 vccd1 _08343_/B sky130_fd_sc_hd__mux2_1
X_05554_ _05076_/A _11428_/Q _11423_/Q _05620_/B2 _05553_/X vssd1 vssd1 vccd1 vccd1
+ _05555_/B sky130_fd_sc_hd__a221o_4
XFILLER_71_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05485_ _10230_/Q input72/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05485_/X sky130_fd_sc_hd__mux2_1
X_08273_ _08793_/A _08273_/B vssd1 vssd1 vccd1 vccd1 _10968_/D sky130_fd_sc_hd__or2_1
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07224_ _07088_/X _10379_/Q _07233_/S vssd1 vssd1 vccd1 vccd1 _10379_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07155_ _07796_/A _07155_/B vssd1 vssd1 vccd1 vccd1 _10338_/D sky130_fd_sc_hd__or2_1
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06106_ _10283_/Q _06106_/B vssd1 vssd1 vccd1 vccd1 _06106_/X sky130_fd_sc_hd__or2_1
XFILLER_69_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07086_ _07664_/A _08645_/S vssd1 vssd1 vccd1 vccd1 _07086_/Y sky130_fd_sc_hd__nor2_4
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06037_ _11806_/Q _06227_/A2 _06035_/X _06036_/X vssd1 vssd1 vccd1 vccd1 _06037_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07988_ _10819_/Q _07991_/S _07363_/S _08817_/B2 vssd1 vssd1 vccd1 vccd1 _10819_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09727_ _11476_/Q _09568_/A _09881_/A2 _11469_/Q vssd1 vssd1 vccd1 vccd1 _09727_/X
+ sky130_fd_sc_hd__a22o_1
X_06939_ _06939_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _08955_/A sky130_fd_sc_hd__or2_2
XFILLER_74_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09658_ _10312_/Q _09566_/B _09571_/D _10315_/Q _09657_/X vssd1 vssd1 vccd1 vccd1
+ _09659_/D sky130_fd_sc_hd__a221o_1
XFILLER_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08609_ _11159_/Q _08633_/B vssd1 vssd1 vccd1 vccd1 _08609_/X sky130_fd_sc_hd__or2_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _10520_/Q _09571_/A _09572_/C _10521_/Q vssd1 vssd1 vccd1 vccd1 _09589_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11620_ _11812_/CLK _11620_/D vssd1 vssd1 vccd1 vccd1 _11620_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11551_ _11763_/CLK _11551_/D vssd1 vssd1 vccd1 vccd1 _11551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10502_ _11439_/CLK _10502_/D vssd1 vssd1 vccd1 vccd1 _10502_/Q sky130_fd_sc_hd__dfxtp_2
X_11482_ _11485_/CLK _11482_/D vssd1 vssd1 vccd1 vccd1 _11482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10433_ _11284_/CLK _10433_/D vssd1 vssd1 vccd1 vccd1 _10433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10364_ _11698_/CLK _10364_/D vssd1 vssd1 vccd1 vccd1 _10364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10295_ _11712_/CLK _10295_/D vssd1 vssd1 vccd1 vccd1 _10295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout690 _11597_/Q vssd1 vssd1 vccd1 vccd1 _05326_/S sky130_fd_sc_hd__buf_12
XFILLER_98_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11749_ _11809_/CLK _11749_/D vssd1 vssd1 vccd1 vccd1 _11749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05270_ _05270_/A _05270_/B vssd1 vssd1 vccd1 vccd1 _05270_/Y sky130_fd_sc_hd__nor2_2
XFILLER_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08960_ _08959_/X _11333_/Q _09830_/B vssd1 vssd1 vccd1 vccd1 _08961_/B sky130_fd_sc_hd__mux2_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07911_ _09129_/A1 _10773_/Q _09206_/B vssd1 vssd1 vccd1 vccd1 _07912_/B sky130_fd_sc_hd__mux2_1
XFILLER_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08891_ _08941_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _11302_/D sky130_fd_sc_hd__or2_1
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07842_ _07042_/A _07819_/Y _07959_/S _10737_/Q vssd1 vssd1 vccd1 vccd1 _10737_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07773_ _10693_/Q _07245_/X _07773_/S vssd1 vssd1 vccd1 vccd1 _10693_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09512_ _09512_/A vssd1 vssd1 vccd1 vccd1 _09512_/Y sky130_fd_sc_hd__inv_2
X_06724_ _10391_/Q _07222_/A _07190_/A _10359_/Q vssd1 vssd1 vccd1 vccd1 _06724_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09443_ input10/X input40/X input17/X input26/X _11576_/Q _11577_/Q vssd1 vssd1 vccd1
+ vccd1 _09443_/X sky130_fd_sc_hd__mux4_1
X_06655_ _06649_/X _06654_/X _11872_/A vssd1 vssd1 vccd1 vccd1 _06655_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05606_ _05630_/A2 _11541_/Q _11538_/Q _05606_/B2 _05604_/X vssd1 vssd1 vccd1 vccd1
+ _05609_/A sky130_fd_sc_hd__a221o_4
X_09374_ _11545_/Q _09376_/B vssd1 vssd1 vccd1 vccd1 _09374_/X sky130_fd_sc_hd__or2_1
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06586_ _10832_/Q _07994_/A _07692_/A _11150_/Q _06585_/X vssd1 vssd1 vccd1 vccd1
+ _06586_/X sky130_fd_sc_hd__o221a_1
XFILLER_71_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08325_ _08439_/A _08325_/B vssd1 vssd1 vccd1 vccd1 _08325_/Y sky130_fd_sc_hd__nand2_4
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05537_ _05537_/A _05537_/B vssd1 vssd1 vccd1 vccd1 _05537_/Y sky130_fd_sc_hd__nor2_8
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08256_ _09283_/A1 _10960_/Q _08276_/S vssd1 vssd1 vccd1 vccd1 _08257_/B sky130_fd_sc_hd__mux2_1
X_05468_ _10757_/Q _09944_/B1 _09872_/B1 _10804_/Q vssd1 vssd1 vccd1 vccd1 _05469_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07207_ _09214_/A _07205_/B _07773_/S _10365_/Q vssd1 vssd1 vccd1 vccd1 _10365_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08187_ _08193_/A _08187_/B vssd1 vssd1 vccd1 vccd1 _10927_/D sky130_fd_sc_hd__or2_1
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05399_ _11220_/Q _11219_/Q _05399_/S vssd1 vssd1 vccd1 vccd1 _05400_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07138_ _10330_/Q _07126_/B _07186_/S _07034_/X vssd1 vssd1 vccd1 vccd1 _10330_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_145_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07069_ _07031_/A _07074_/S _07068_/X _07141_/B vssd1 vssd1 vccd1 vccd1 _10293_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10080_ _10080_/A0 _11740_/Q _10082_/S vssd1 vssd1 vccd1 vccd1 _11740_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10982_ _11307_/CLK _10982_/D vssd1 vssd1 vccd1 vccd1 _10982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11603_ _11604_/CLK _11603_/D vssd1 vssd1 vccd1 vccd1 _11603_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11534_ _11762_/CLK _11534_/D vssd1 vssd1 vccd1 vccd1 _11534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11465_ _11465_/CLK _11465_/D vssd1 vssd1 vccd1 vccd1 _11465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10416_ _11439_/CLK _10416_/D vssd1 vssd1 vccd1 vccd1 _10416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11396_ _11410_/CLK _11396_/D vssd1 vssd1 vccd1 vccd1 _11396_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10347_ _11465_/CLK _10347_/D vssd1 vssd1 vccd1 vccd1 _10347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10278_ _11474_/CLK _10278_/D vssd1 vssd1 vccd1 vccd1 _10278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06440_ _10484_/Q _08649_/A _06437_/X _06439_/X vssd1 vssd1 vccd1 vccd1 _06440_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06371_ _10623_/Q _06371_/A2 _06998_/A _10510_/Q vssd1 vssd1 vccd1 vccd1 _06374_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08110_ _10880_/Q _08120_/S _07642_/S _08811_/B2 vssd1 vssd1 vccd1 vccd1 _10880_/D
+ sky130_fd_sc_hd__o22a_1
X_05322_ _10882_/Q _10881_/Q _05394_/S vssd1 vssd1 vccd1 vccd1 _05323_/D sky130_fd_sc_hd__mux2_1
X_09090_ _09090_/A1 _09082_/X _09089_/X _09092_/C1 vssd1 vssd1 vccd1 vccd1 _11392_/D
+ sky130_fd_sc_hd__o211a_1
X_08041_ _10845_/Q _08051_/S _07365_/Y _07232_/B vssd1 vssd1 vccd1 vccd1 _10845_/D
+ sky130_fd_sc_hd__o22a_1
X_05253_ _05253_/A _05253_/B _05253_/C _05253_/D vssd1 vssd1 vccd1 vccd1 _05259_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_31_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05184_ _05184_/A _05184_/B _05184_/C _05184_/D vssd1 vssd1 vccd1 vccd1 _05190_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_143_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09992_ _11683_/Q _09994_/B vssd1 vssd1 vccd1 vccd1 _09992_/X sky130_fd_sc_hd__or2_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08943_ _09237_/A0 _08940_/S _08942_/X _08943_/C1 vssd1 vssd1 vccd1 vccd1 _11330_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08874_ _09101_/A1 _11294_/Q _08874_/S vssd1 vssd1 vccd1 vccd1 _08875_/B sky130_fd_sc_hd__mux2_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07825_ _10021_/A0 _07839_/A2 _07961_/S _10720_/Q vssd1 vssd1 vccd1 vccd1 _10720_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07756_ _10679_/Q _07760_/B vssd1 vssd1 vccd1 vccd1 _07756_/X sky130_fd_sc_hd__or2_1
XFILLER_129_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06707_ _10572_/Q _06806_/A2 _06728_/B1 _10501_/Q _06706_/X vssd1 vssd1 vccd1 vccd1
+ _06707_/X sky130_fd_sc_hd__o221a_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07687_ _10643_/Q _07673_/Y _07676_/X _07316_/X vssd1 vssd1 vccd1 vccd1 _10643_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09426_ _11642_/Q _11585_/Q _09426_/S vssd1 vssd1 vccd1 vccd1 _11585_/D sky130_fd_sc_hd__mux2_1
X_06638_ _11180_/Q _08647_/B _06634_/X _06637_/X vssd1 vssd1 vccd1 vccd1 _06644_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09357_ _10118_/A0 _11537_/Q _09357_/S vssd1 vssd1 vccd1 vccd1 _11537_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06569_ _06560_/X _06563_/X _06568_/X vssd1 vssd1 vccd1 vccd1 _06569_/X sky130_fd_sc_hd__o21a_2
XFILLER_21_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08308_ _10988_/Q _08301_/Y _08304_/Y _07227_/X vssd1 vssd1 vccd1 vccd1 _10988_/D
+ sky130_fd_sc_hd__a22o_1
X_09288_ _11496_/Q _09288_/B vssd1 vssd1 vccd1 vccd1 _09288_/X sky130_fd_sc_hd__or2_1
XFILLER_100_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08239_ _08760_/A0 _10953_/Q _08325_/B vssd1 vssd1 vccd1 vccd1 _08240_/B sky130_fd_sc_hd__mux2_1
XFILLER_153_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11250_ _11428_/CLK _11250_/D vssd1 vssd1 vccd1 vccd1 _11250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10201_ _11803_/CLK _10201_/D vssd1 vssd1 vccd1 vccd1 _10201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11181_ _11307_/CLK _11181_/D vssd1 vssd1 vccd1 vccd1 _11181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10132_ _10132_/A0 _11778_/Q _10135_/S vssd1 vssd1 vccd1 vccd1 _11778_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10063_ _10110_/A0 _11724_/Q _10071_/S vssd1 vssd1 vccd1 vccd1 _11724_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10965_ _11572_/CLK _10965_/D vssd1 vssd1 vccd1 vccd1 _10965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10896_ _11632_/CLK _10896_/D vssd1 vssd1 vccd1 vccd1 _10896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11517_ _11756_/CLK _11517_/D vssd1 vssd1 vccd1 vccd1 _11517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11448_ _11450_/CLK _11448_/D vssd1 vssd1 vccd1 vccd1 _11448_/Q sky130_fd_sc_hd__dfxtp_1
X_11379_ _11428_/CLK _11379_/D vssd1 vssd1 vccd1 vccd1 _11379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05940_ _10822_/Q _06415_/A2 _06628_/B1 _10987_/Q vssd1 vssd1 vccd1 vccd1 _05940_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05871_ _10418_/Q _06318_/A2 _06504_/B1 _11001_/Q vssd1 vssd1 vccd1 vccd1 _05871_/X
+ sky130_fd_sc_hd__o22a_1
X_07610_ _10590_/Q _07598_/Y _07599_/Y _07318_/X vssd1 vssd1 vccd1 vccd1 _10590_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08590_ _08590_/A _08590_/B vssd1 vssd1 vccd1 vccd1 _11150_/D sky130_fd_sc_hd__or2_1
XFILLER_94_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07541_ _07303_/A _10554_/Q _07589_/S vssd1 vssd1 vccd1 vccd1 _07542_/B sky130_fd_sc_hd__mux2_1
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07472_ input92/X _10514_/Q _07477_/S vssd1 vssd1 vccd1 vccd1 _07473_/B sky130_fd_sc_hd__mux2_1
X_09211_ _11453_/Q _09206_/Y _09208_/Y _07013_/X vssd1 vssd1 vccd1 vccd1 _11453_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06423_ _10739_/Q _07202_/A _05865_/B _11776_/Q _06422_/X vssd1 vssd1 vccd1 vccd1
+ _06423_/X sky130_fd_sc_hd__o221a_1
XFILLER_50_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09142_ _11416_/Q _09132_/X _09141_/X vssd1 vssd1 vccd1 vccd1 _11416_/D sky130_fd_sc_hd__a21o_1
X_06354_ _11398_/Q _06716_/A2 _09110_/A _11411_/Q vssd1 vssd1 vccd1 vccd1 _06354_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_72_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05305_ _11014_/Q _11013_/Q _11595_/Q vssd1 vssd1 vccd1 vccd1 _05307_/C sky130_fd_sc_hd__mux2_1
XFILLER_135_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09073_ _11385_/Q _09077_/B vssd1 vssd1 vccd1 vccd1 _09073_/X sky130_fd_sc_hd__or2_1
XFILLER_120_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06285_ _11367_/Q _09016_/A _08994_/A _11357_/Q _07689_/B vssd1 vssd1 vccd1 vccd1
+ _06285_/X sky130_fd_sc_hd__o221a_1
X_08024_ _09141_/A1 _08035_/S _08023_/X _08791_/C1 vssd1 vssd1 vccd1 vccd1 _10836_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05236_ _05419_/S _11009_/Q _11008_/Q _09679_/B _05230_/X vssd1 vssd1 vccd1 vccd1
+ _05238_/C sky130_fd_sc_hd__a221oi_2
XFILLER_151_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05167_ _05167_/A _05167_/B _05167_/C _05167_/D vssd1 vssd1 vccd1 vccd1 _05168_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_103_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09975_ _10190_/A0 _11675_/Q _09975_/S vssd1 vssd1 vccd1 vccd1 _11675_/D sky130_fd_sc_hd__mux2_1
X_05098_ _11576_/Q vssd1 vssd1 vccd1 vccd1 _09441_/A sky130_fd_sc_hd__inv_2
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08926_ _11322_/Q _08946_/B vssd1 vssd1 vccd1 vccd1 _08926_/X sky130_fd_sc_hd__or2_1
XFILLER_103_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08857_ _08869_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _11285_/D sky130_fd_sc_hd__or2_1
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07808_ _07930_/A _07808_/B vssd1 vssd1 vccd1 vccd1 _10711_/D sky130_fd_sc_hd__or2_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _11250_/Q _08804_/B vssd1 vssd1 vccd1 vccd1 _08788_/X sky130_fd_sc_hd__or2_1
XFILLER_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ _07028_/A _07761_/A2 _07738_/X _09201_/A1 vssd1 vssd1 vccd1 vccd1 _10670_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _11622_/CLK _10750_/D vssd1 vssd1 vccd1 vccd1 _10750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09409_ _11654_/Q _11570_/Q _09414_/S vssd1 vssd1 vccd1 vccd1 _11570_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10681_ _11457_/CLK _10681_/D vssd1 vssd1 vccd1 vccd1 _10681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_wb_clk_i clkbuf_leaf_69_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11792_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11302_ _11330_/CLK _11302_/D vssd1 vssd1 vccd1 vccd1 _11302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11233_ _11233_/CLK _11233_/D vssd1 vssd1 vccd1 vccd1 _11233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11164_ _11243_/CLK _11164_/D vssd1 vssd1 vccd1 vccd1 _11164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10115_ _10115_/A0 _11762_/Q _10118_/S vssd1 vssd1 vccd1 vccd1 _11762_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11095_ _11675_/CLK _11095_/D vssd1 vssd1 vccd1 vccd1 _11095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10046_ _10050_/A _10046_/B vssd1 vssd1 vccd1 vccd1 _11714_/D sky130_fd_sc_hd__or2_1
XFILLER_76_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10948_ _11023_/CLK _10948_/D vssd1 vssd1 vccd1 vccd1 _10948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10879_ _10929_/CLK _10879_/D vssd1 vssd1 vccd1 vccd1 _10879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _05224_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06070_ _10824_/Q _07994_/A _08300_/A _11269_/Q vssd1 vssd1 vccd1 vccd1 _06070_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout508 _09048_/C1 vssd1 vssd1 vccd1 vccd1 _09279_/C1 sky130_fd_sc_hd__clkbuf_8
Xfanout519 _07420_/A vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__buf_8
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09760_ input6/X _09740_/Y _09759_/X vssd1 vssd1 vccd1 vccd1 _09760_/X sky130_fd_sc_hd__a21o_1
XFILLER_100_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ _06970_/X _06971_/Y _06950_/A vssd1 vssd1 vccd1 vccd1 _06972_/X sky130_fd_sc_hd__o21a_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _11210_/Q _08718_/S _07852_/S _07227_/B vssd1 vssd1 vccd1 vccd1 _11210_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05923_ _11191_/Q _09154_/A _08594_/A _11154_/Q _05922_/X vssd1 vssd1 vccd1 vccd1
+ _05923_/X sky130_fd_sc_hd__o221a_2
X_09691_ _09703_/A _09691_/B vssd1 vssd1 vccd1 vccd1 _11637_/D sky130_fd_sc_hd__or2_1
XFILLER_6_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08642_ _11176_/Q _08645_/S _07086_/Y _07227_/B vssd1 vssd1 vccd1 vccd1 _11176_/D
+ sky130_fd_sc_hd__o22a_1
X_05854_ _05851_/X _05852_/X _05853_/X _05848_/X vssd1 vssd1 vccd1 vccd1 _05854_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _08745_/A _08573_/B vssd1 vssd1 vccd1 vccd1 _11141_/D sky130_fd_sc_hd__or2_1
X_05785_ _05779_/X _05784_/X _07151_/B vssd1 vssd1 vccd1 vccd1 _05785_/X sky130_fd_sc_hd__o21a_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07524_ _07922_/A _07524_/B vssd1 vssd1 vccd1 vccd1 _10546_/D sky130_fd_sc_hd__or2_1
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07455_ _07455_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07455_/X sky130_fd_sc_hd__or2_4
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06406_ _06663_/A _10231_/Q vssd1 vssd1 vccd1 vccd1 _06406_/X sky130_fd_sc_hd__and2_1
X_07386_ _08749_/A _07386_/B vssd1 vssd1 vccd1 vccd1 _10468_/D sky130_fd_sc_hd__or2_1
X_09125_ _10023_/A0 _09127_/B _09129_/B1 vssd1 vssd1 vccd1 vccd1 _09125_/X sky130_fd_sc_hd__a21o_1
X_06337_ _06328_/X _06331_/X _06336_/X vssd1 vssd1 vccd1 vccd1 _06337_/X sky130_fd_sc_hd__a21o_2
XFILLER_136_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09056_ _09172_/A1 _09038_/X _09055_/X _09289_/C1 vssd1 vssd1 vccd1 vccd1 _11377_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06268_ _11060_/Q _06631_/A2 _06632_/A2 _11174_/Q _06392_/C1 vssd1 vssd1 vccd1 vccd1
+ _06268_/X sky130_fd_sc_hd__o221a_1
X_08007_ _10828_/Q _08091_/C vssd1 vssd1 vccd1 vccd1 _08007_/X sky130_fd_sc_hd__or2_1
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05219_ _06941_/A _10860_/Q _10853_/Q _05377_/S vssd1 vssd1 vccd1 vccd1 _05224_/B
+ sky130_fd_sc_hd__a22o_2
X_06199_ _10269_/Q _06999_/A _06195_/X _06198_/X vssd1 vssd1 vccd1 vccd1 _06199_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09958_ _09958_/A _09958_/B vssd1 vssd1 vccd1 vccd1 _09959_/C sky130_fd_sc_hd__nor2_4
XFILLER_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ _09111_/A1 _08945_/A2 _08908_/X _08919_/C1 vssd1 vssd1 vccd1 vccd1 _11313_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_114_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11712_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09889_ _09889_/A vssd1 vssd1 vccd1 vccd1 _09889_/Y sky130_fd_sc_hd__clkinv_2
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_tms1x00_1100 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1100/HI io_oeb[30] sky130_fd_sc_hd__conb_1
XFILLER_131_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_tms1x00_1111 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1111/HI io_out[3] sky130_fd_sc_hd__conb_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1122 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1122/HI irq[2] sky130_fd_sc_hd__conb_1
XFILLER_73_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _11720_/CLK _10802_/D vssd1 vssd1 vccd1 vccd1 _10802_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _11791_/CLK _11782_/D vssd1 vssd1 vccd1 vccd1 _11782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10733_ _11722_/CLK _10733_/D vssd1 vssd1 vccd1 vccd1 _10733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10664_ _11644_/CLK _10664_/D vssd1 vssd1 vccd1 vccd1 _10664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10595_ _11243_/CLK _10595_/D vssd1 vssd1 vccd1 vccd1 _10595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11216_ _11220_/CLK _11216_/D vssd1 vssd1 vccd1 vccd1 _11216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ _11151_/CLK _11147_/D vssd1 vssd1 vccd1 vccd1 _11147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11078_ _11766_/CLK _11078_/D vssd1 vssd1 vccd1 vccd1 _11078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10029_ _11704_/Q _10051_/S _10027_/Y _07314_/B vssd1 vssd1 vccd1 vccd1 _11704_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05570_ _05616_/A1 _11419_/Q _11416_/Q _05077_/A _05569_/X vssd1 vssd1 vccd1 vccd1
+ _05573_/A sky130_fd_sc_hd__a221o_4
XFILLER_32_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07240_ _10388_/Q _07233_/S _07239_/X _09206_/A vssd1 vssd1 vccd1 vccd1 _10388_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07171_ _07934_/A _07171_/B vssd1 vssd1 vccd1 vccd1 _10346_/D sky130_fd_sc_hd__or2_1
X_06122_ _10878_/Q _06513_/A2 _06636_/A2 _10926_/Q _07083_/B vssd1 vssd1 vccd1 vccd1
+ _06125_/B sky130_fd_sc_hd__o221a_2
XFILLER_121_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06053_ _11156_/Q _08594_/A _06718_/C1 _06052_/X vssd1 vssd1 vccd1 vccd1 _06053_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout305 _07540_/X vssd1 vssd1 vccd1 vccd1 _07557_/S sky130_fd_sc_hd__buf_6
XFILLER_67_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout316 _07364_/X vssd1 vssd1 vccd1 vccd1 _08051_/S sky130_fd_sc_hd__buf_6
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout327 _07425_/S vssd1 vssd1 vccd1 vccd1 _07429_/S sky130_fd_sc_hd__buf_8
X_09812_ _10297_/Q _09571_/A _09573_/D _10284_/Q vssd1 vssd1 vccd1 vccd1 _09815_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout338 _07483_/S vssd1 vssd1 vccd1 vccd1 _07477_/S sky130_fd_sc_hd__buf_8
XFILLER_115_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout349 _08230_/B vssd1 vssd1 vccd1 vccd1 _08665_/C sky130_fd_sc_hd__buf_8
XFILLER_115_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09743_ _10498_/Q _09886_/A2 _09872_/B1 _10535_/Q vssd1 vssd1 vccd1 vccd1 _09743_/X
+ sky130_fd_sc_hd__a22o_1
X_06955_ _08956_/B _06954_/X _06969_/S vssd1 vssd1 vccd1 vccd1 _06955_/X sky130_fd_sc_hd__mux2_4
XFILLER_132_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05906_ _05903_/X _05905_/X _05901_/X vssd1 vssd1 vccd1 vccd1 _05906_/X sky130_fd_sc_hd__a21o_2
X_09674_ _09674_/A vssd1 vssd1 vccd1 vccd1 _09674_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06886_ _07092_/A _06886_/A2 _06884_/Y _10216_/Q vssd1 vssd1 vccd1 vccd1 _10216_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08625_ _11167_/Q _08633_/B vssd1 vssd1 vccd1 vccd1 _08625_/X sky130_fd_sc_hd__or2_1
X_05837_ _11559_/Q _09391_/A _06284_/B1 _11549_/Q vssd1 vssd1 vccd1 vccd1 _05837_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08556_ _11132_/Q _08558_/S _07355_/S _07316_/B vssd1 vssd1 vccd1 vccd1 _11132_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05768_ _11558_/Q _09391_/A _09380_/A _11548_/Q vssd1 vssd1 vccd1 vccd1 _05768_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07507_ _10538_/Q _07537_/B vssd1 vssd1 vccd1 vccd1 _07507_/X sky130_fd_sc_hd__or2_1
XFILLER_35_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08487_ _10080_/A0 _11094_/Q _08497_/S vssd1 vssd1 vccd1 vccd1 _08488_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05699_ _11105_/Q _05531_/Y _05567_/Y _11106_/Q vssd1 vssd1 vccd1 vccd1 _05699_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07438_ _10058_/A _07438_/B vssd1 vssd1 vccd1 vccd1 _10495_/D sky130_fd_sc_hd__or2_1
XFILLER_91_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07369_ _10457_/Q _07090_/X _07373_/S vssd1 vssd1 vccd1 vccd1 _10457_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09108_ _07043_/B _07539_/Y _09107_/X vssd1 vssd1 vccd1 vccd1 _11401_/D sky130_fd_sc_hd__a21o_1
X_10380_ _10981_/CLK _10380_/D vssd1 vssd1 vccd1 vccd1 _10380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ _09111_/A1 _09055_/B _09290_/B1 vssd1 vssd1 vccd1 vccd1 _09039_/X sky130_fd_sc_hd__a21o_1
XFILLER_2_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11001_ _11005_/CLK _11001_/D vssd1 vssd1 vccd1 vccd1 _11001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout850 fanout861/X vssd1 vssd1 vccd1 vccd1 _06635_/A2 sky130_fd_sc_hd__buf_6
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout861 _05741_/Y vssd1 vssd1 vccd1 vccd1 fanout861/X sky130_fd_sc_hd__buf_8
Xfanout872 _06719_/A2 vssd1 vssd1 vccd1 vccd1 _06736_/A2 sky130_fd_sc_hd__buf_6
Xfanout883 _06227_/A2 vssd1 vssd1 vccd1 vccd1 _06631_/A2 sky130_fd_sc_hd__buf_4
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout894 _06539_/A2 vssd1 vssd1 vccd1 vccd1 _06454_/A2 sky130_fd_sc_hd__buf_4
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _11765_/CLK _11765_/D vssd1 vssd1 vccd1 vccd1 _11765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_82_wb_clk_i clkbuf_leaf_85_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11575_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _10765_/CLK _10716_/D vssd1 vssd1 vccd1 vccd1 _10716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11696_ _11713_/CLK _11696_/D vssd1 vssd1 vccd1 vccd1 _11696_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11629_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ _11270_/CLK _10647_/D vssd1 vssd1 vccd1 vccd1 _10647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10578_ _10765_/CLK _10578_/D vssd1 vssd1 vccd1 vccd1 _10578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06740_ _06577_/A _10241_/Q _06855_/B vssd1 vssd1 vccd1 vccd1 _06740_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06671_ _11444_/Q _07778_/A _06727_/B _10407_/Q vssd1 vssd1 vccd1 vccd1 _06671_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08410_ _11046_/Q _08422_/B vssd1 vssd1 vccd1 vccd1 _08410_/X sky130_fd_sc_hd__or2_1
X_05622_ _11753_/Q _05628_/A2 _05628_/B1 _11750_/Q vssd1 vssd1 vccd1 vccd1 _05622_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09390_ _10118_/A0 _11557_/Q _09390_/S vssd1 vssd1 vccd1 vccd1 _11557_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08341_ _08579_/A0 _08360_/S _08340_/X _09022_/C1 vssd1 vssd1 vccd1 vccd1 _11013_/D
+ sky130_fd_sc_hd__o211a_1
X_05553_ _05619_/A1 _11431_/Q _11427_/Q _05619_/B2 _05551_/X vssd1 vssd1 vccd1 vccd1
+ _05553_/X sky130_fd_sc_hd__a221o_1
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08272_ _08935_/A1 _10968_/Q _08272_/S vssd1 vssd1 vccd1 vccd1 _08273_/B sky130_fd_sc_hd__mux2_1
X_05484_ _10229_/Q input71/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05484_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07223_ _07664_/A _07663_/S vssd1 vssd1 vccd1 vccd1 _07223_/Y sky130_fd_sc_hd__nor2_2
XFILLER_121_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07154_ _07303_/A _10338_/Q _07172_/S vssd1 vssd1 vccd1 vccd1 _07155_/B sky130_fd_sc_hd__mux2_1
XFILLER_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06105_ _10621_/Q _06371_/A2 _06105_/B1 _10797_/Q vssd1 vssd1 vccd1 vccd1 _06105_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_156_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07085_ _08286_/A _08560_/C _07847_/C vssd1 vssd1 vccd1 vccd1 _08645_/S sky130_fd_sc_hd__and3_4
XFILLER_106_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06036_ _10260_/Q _06976_/A _06903_/A _10197_/Q vssd1 vssd1 vccd1 vccd1 _06036_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07987_ _08196_/A _07987_/B vssd1 vssd1 vccd1 vccd1 _10818_/D sky130_fd_sc_hd__or2_1
XFILLER_87_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09726_ _10351_/Q _09878_/A2 _09872_/B1 _11464_/Q _09725_/X vssd1 vssd1 vccd1 vccd1
+ _09731_/B sky130_fd_sc_hd__a221o_1
X_06938_ _09703_/A _06938_/B vssd1 vssd1 vccd1 vccd1 _09416_/A sky130_fd_sc_hd__nor2_8
XFILLER_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09657_ _10320_/Q _09947_/A2 _09568_/B _10314_/Q vssd1 vssd1 vccd1 vccd1 _09657_/X
+ sky130_fd_sc_hd__a22o_1
X_06869_ _10337_/Q _07539_/A vssd1 vssd1 vccd1 vccd1 _06869_/X sky130_fd_sc_hd__or2_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _08682_/A _08608_/B vssd1 vssd1 vccd1 vccd1 _11158_/D sky130_fd_sc_hd__or2_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _10275_/Q _09567_/B _09947_/B1 _10516_/Q _09587_/X vssd1 vssd1 vccd1 vccd1
+ _09593_/A sky130_fd_sc_hd__a221o_1
XFILLER_63_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _11119_/Q _08545_/B vssd1 vssd1 vccd1 vccd1 _08539_/X sky130_fd_sc_hd__or2_1
XFILLER_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11550_ _11758_/CLK _11550_/D vssd1 vssd1 vccd1 vccd1 _11550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ _11470_/CLK _10501_/D vssd1 vssd1 vccd1 vccd1 _10501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11481_ _11485_/CLK _11481_/D vssd1 vssd1 vccd1 vccd1 _11481_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10432_ _11284_/CLK _10432_/D vssd1 vssd1 vccd1 vccd1 _10432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10363_ _11745_/CLK _10363_/D vssd1 vssd1 vccd1 vccd1 _10363_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_100_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10294_ _10725_/CLK _10294_/D vssd1 vssd1 vccd1 vccd1 _10294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout680 _11599_/Q vssd1 vssd1 vccd1 vccd1 _05413_/S sky130_fd_sc_hd__buf_12
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout691 _05372_/S vssd1 vssd1 vccd1 vccd1 _05393_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _11755_/CLK _11748_/D vssd1 vssd1 vccd1 vccd1 _11748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11679_ _11684_/CLK _11679_/D vssd1 vssd1 vccd1 vccd1 _11679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07910_ _07928_/A _07910_/B vssd1 vssd1 vccd1 vccd1 _10772_/D sky130_fd_sc_hd__or2_1
XFILLER_68_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08890_ _09237_/A0 _11302_/Q _08890_/S vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07841_ _07147_/A _07819_/Y _07961_/S _10736_/Q vssd1 vssd1 vccd1 vccd1 _10736_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07772_ _10692_/Q _07241_/X _07772_/S vssd1 vssd1 vccd1 vccd1 _10692_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06723_ _06704_/B _06722_/X _06704_/Y vssd1 vssd1 vccd1 vccd1 _10240_/D sky130_fd_sc_hd__o21ai_1
X_09511_ _09515_/C _09515_/B _09511_/C vssd1 vssd1 vccd1 vccd1 _09512_/A sky130_fd_sc_hd__and3b_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09442_ _11576_/Q _11577_/Q vssd1 vssd1 vccd1 vccd1 _09442_/X sky130_fd_sc_hd__or2_2
X_06654_ _11710_/Q _08560_/A _06650_/X _06653_/X vssd1 vssd1 vccd1 vccd1 _06654_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05605_ _05629_/A2 _11546_/Q _11540_/Q _05629_/B1 vssd1 vssd1 vccd1 vccd1 _05605_/X
+ sky130_fd_sc_hd__a22o_1
X_09373_ _11544_/Q _09359_/X _09372_/X vssd1 vssd1 vccd1 vccd1 _11544_/D sky130_fd_sc_hd__a21o_1
XFILLER_36_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06585_ _10859_/Q _08054_/A vssd1 vssd1 vccd1 vccd1 _06585_/X sky130_fd_sc_hd__or2_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08324_ _08438_/A _08324_/B vssd1 vssd1 vccd1 vccd1 _08324_/Y sky130_fd_sc_hd__nor2_1
X_05536_ _05626_/A2 _11524_/Q _11519_/Q _05630_/B1 _05535_/X vssd1 vssd1 vccd1 vccd1
+ _05537_/B sky130_fd_sc_hd__a221o_4
XFILLER_71_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08255_ _08851_/A _08255_/B vssd1 vssd1 vccd1 vccd1 _10959_/D sky130_fd_sc_hd__or2_1
X_05467_ _10808_/Q _09572_/B _09878_/A2 _10763_/Q _05459_/X vssd1 vssd1 vccd1 vccd1
+ _05469_/C sky130_fd_sc_hd__a221o_1
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07206_ _07303_/A _07205_/B _07773_/S _10364_/Q vssd1 vssd1 vccd1 vccd1 _10364_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08186_ _10927_/Q _07015_/A _08197_/S vssd1 vssd1 vccd1 vccd1 _08187_/B sky130_fd_sc_hd__mux2_1
XFILLER_118_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05398_ _10745_/Q _10744_/Q _05398_/S vssd1 vssd1 vccd1 vccd1 _05400_/C sky130_fd_sc_hd__mux2_1
XFILLER_134_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07137_ _10047_/A1 _07111_/X _07136_/X _07147_/B vssd1 vssd1 vccd1 vccd1 _10329_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07068_ _10293_/Q _07078_/B vssd1 vssd1 vccd1 vccd1 _07068_/X sky130_fd_sc_hd__or2_1
XFILLER_47_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06019_ _11750_/Q _10087_/A _10137_/A _11786_/Q _06214_/C1 vssd1 vssd1 vccd1 vccd1
+ _06019_/X sky130_fd_sc_hd__o221a_2
XFILLER_102_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09709_ _11434_/Q _09877_/A2 _09573_/A _10404_/Q vssd1 vssd1 vccd1 vccd1 _09709_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_90_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10981_ _10981_/CLK _10981_/D vssd1 vssd1 vccd1 vccd1 _10981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11602_ _11604_/CLK _11602_/D vssd1 vssd1 vccd1 vccd1 _11602_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_70_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11533_ _11762_/CLK _11533_/D vssd1 vssd1 vccd1 vccd1 _11533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11464_ _11465_/CLK _11464_/D vssd1 vssd1 vccd1 vccd1 _11464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10415_ _11457_/CLK _10415_/D vssd1 vssd1 vccd1 vccd1 _10415_/Q sky130_fd_sc_hd__dfxtp_1
X_11395_ _11411_/CLK _11395_/D vssd1 vssd1 vccd1 vccd1 _11395_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10346_ _10769_/CLK _10346_/D vssd1 vssd1 vccd1 vccd1 _10346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10277_ _11722_/CLK _10277_/D vssd1 vssd1 vccd1 vccd1 _10277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06370_ _10366_/Q _06370_/A2 _07827_/A2 _10722_/Q vssd1 vssd1 vccd1 vccd1 _06370_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05321_ _10887_/Q _10886_/Q _05399_/S vssd1 vssd1 vccd1 vccd1 _05323_/C sky130_fd_sc_hd__mux2_1
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ _08733_/A _08040_/B vssd1 vssd1 vccd1 vccd1 _10844_/D sky130_fd_sc_hd__or2_1
XFILLER_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05252_ _11082_/Q _11081_/Q _05377_/S vssd1 vssd1 vccd1 vccd1 _05253_/D sky130_fd_sc_hd__mux2_2
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05183_ _10593_/Q _10836_/Q _08956_/B vssd1 vssd1 vccd1 vccd1 _05184_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09991_ _11682_/Q _09977_/X _09990_/X vssd1 vssd1 vccd1 vccd1 _11682_/D sky130_fd_sc_hd__a21o_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08942_ _11330_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08942_/X sky130_fd_sc_hd__or2_1
XFILLER_130_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08873_ _08873_/A _08873_/B vssd1 vssd1 vccd1 vccd1 _11293_/D sky130_fd_sc_hd__or2_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07824_ _07092_/A _07820_/B _07821_/A _10719_/Q vssd1 vssd1 vccd1 vccd1 _10719_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07755_ _07143_/A _07755_/A2 _07754_/X _07868_/C1 vssd1 vssd1 vccd1 vccd1 _10678_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06706_ _10760_/Q _06861_/B _06806_/B1 _10671_/Q vssd1 vssd1 vccd1 vccd1 _06706_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_71_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07686_ _10642_/Q _07674_/X _07675_/Y _07314_/X vssd1 vssd1 vccd1 vccd1 _10642_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06637_ _11220_/Q _06637_/A2 _06636_/X _11869_/A vssd1 vssd1 vccd1 vccd1 _06637_/X
+ sky130_fd_sc_hd__o211a_1
X_09425_ _11641_/Q _11584_/Q _09704_/B vssd1 vssd1 vccd1 vccd1 _11584_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09356_ _10117_/A0 _11536_/Q _09357_/S vssd1 vssd1 vccd1 vccd1 _11536_/D sky130_fd_sc_hd__mux2_1
X_06568_ _10357_/Q _08649_/A _06564_/X _06567_/X vssd1 vssd1 vccd1 vccd1 _06568_/X
+ sky130_fd_sc_hd__a211o_4
Xclkbuf_leaf_139_wb_clk_i clkbuf_4_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11768_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_05519_ _05616_/A1 _11409_/Q _11406_/Q _05077_/A vssd1 vssd1 vccd1 vccd1 _05519_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08307_ _10987_/Q _08302_/Y _08303_/Y _07090_/X vssd1 vssd1 vccd1 vccd1 _10987_/D
+ sky130_fd_sc_hd__o22a_1
X_09287_ _11495_/Q _09271_/X _09286_/X vssd1 vssd1 vccd1 vccd1 _11495_/D sky130_fd_sc_hd__a21o_1
XFILLER_21_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06499_ _10897_/Q _06632_/A2 _06497_/X _06498_/X vssd1 vssd1 vccd1 vccd1 _06499_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08238_ _10150_/A1 _08325_/B _08237_/X _08753_/C1 vssd1 vssd1 vccd1 vccd1 _10952_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08169_ _07007_/A _10911_/Q _08182_/S vssd1 vssd1 vccd1 vccd1 _10911_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10200_ _11803_/CLK _10200_/D vssd1 vssd1 vccd1 vccd1 _10200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11180_ _11268_/CLK _11180_/D vssd1 vssd1 vccd1 vccd1 _11180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10131_ _07061_/A _11777_/Q _10135_/S vssd1 vssd1 vccd1 vccd1 _11777_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10062_ _10181_/A0 _11723_/Q _10071_/S vssd1 vssd1 vccd1 vccd1 _11723_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10964_ _11572_/CLK _10964_/D vssd1 vssd1 vccd1 vccd1 _10964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10895_ _11632_/CLK _10895_/D vssd1 vssd1 vccd1 vccd1 _10895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11516_ _11763_/CLK _11516_/D vssd1 vssd1 vccd1 vccd1 _11516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11447_ _11458_/CLK _11447_/D vssd1 vssd1 vccd1 vccd1 _11447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11378_ _11431_/CLK _11378_/D vssd1 vssd1 vccd1 vccd1 _11378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10329_ _11719_/CLK _10329_/D vssd1 vssd1 vccd1 vccd1 _10329_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05870_ _05866_/X _05869_/X _07083_/A _05864_/X vssd1 vssd1 vccd1 vccd1 _05870_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07540_ _07540_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07540_/X sky130_fd_sc_hd__or2_1
X_07471_ _10513_/Q _07000_/B _07000_/Y _07333_/B vssd1 vssd1 vccd1 vccd1 _10513_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06422_ _11132_/Q _06635_/A2 _06514_/A2 _10605_/Q vssd1 vssd1 vccd1 vccd1 _06422_/X
+ sky130_fd_sc_hd__o22a_1
X_09210_ _11452_/Q _09205_/Y _09209_/Y _07005_/X vssd1 vssd1 vccd1 vccd1 _11452_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09141_ _09141_/A1 _09149_/B _10166_/B1 vssd1 vssd1 vccd1 vccd1 _09141_/X sky130_fd_sc_hd__a21o_1
X_06353_ _07690_/A _06353_/B _06353_/C vssd1 vssd1 vccd1 vccd1 _06353_/X sky130_fd_sc_hd__or3_4
XFILLER_37_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05304_ _10874_/Q _10873_/Q _05326_/S vssd1 vssd1 vccd1 vccd1 _05307_/B sky130_fd_sc_hd__mux2_1
X_09072_ _11384_/Q _09060_/X _09071_/X vssd1 vssd1 vccd1 vccd1 _11384_/D sky130_fd_sc_hd__a21o_1
X_06284_ _11566_/Q _09391_/A _06284_/B1 _11556_/Q _06283_/X vssd1 vssd1 vccd1 vccd1
+ _06284_/X sky130_fd_sc_hd__o221a_1
XFILLER_129_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08023_ _10836_/Q _08037_/B vssd1 vssd1 vccd1 vccd1 _08023_/X sky130_fd_sc_hd__or2_1
X_05235_ _05471_/A _08241_/A _05231_/Y _05232_/Y _05234_/Y vssd1 vssd1 vccd1 vccd1
+ _05238_/B sky130_fd_sc_hd__o2111a_1
XFILLER_116_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05166_ _11078_/Q _10598_/Q _05385_/S vssd1 vssd1 vccd1 vccd1 _05167_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09974_ _10117_/A0 _11674_/Q _09975_/S vssd1 vssd1 vccd1 vccd1 _11674_/D sky130_fd_sc_hd__mux2_1
X_05097_ _09540_/A vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__clkinv_4
XFILLER_104_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08925_ _09172_/A1 _08940_/S _08924_/X _09122_/C1 vssd1 vssd1 vccd1 vccd1 _11321_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08856_ _09111_/A1 _11285_/Q _08874_/S vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__mux2_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07807_ _08423_/A1 _10711_/Q _09193_/B vssd1 vssd1 vccd1 vccd1 _07808_/B sky130_fd_sc_hd__mux2_1
XFILLER_57_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05999_ _10604_/Q _06635_/B1 _05995_/X _05998_/X vssd1 vssd1 vccd1 vccd1 _06000_/C
+ sky130_fd_sc_hd__o211a_2
X_08787_ _08875_/A _08787_/B vssd1 vssd1 vccd1 vccd1 _11249_/D sky130_fd_sc_hd__or2_1
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ _10670_/Q _07760_/B vssd1 vssd1 vccd1 vccd1 _07738_/X sky130_fd_sc_hd__or2_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07669_ _10630_/Q _07665_/S _07249_/S _07451_/B vssd1 vssd1 vccd1 vccd1 _10630_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09408_ _11653_/Q _11569_/Q _09414_/S vssd1 vssd1 vccd1 vccd1 _11569_/D sky130_fd_sc_hd__mux2_1
X_10680_ _11439_/CLK _10680_/D vssd1 vssd1 vccd1 vccd1 _10680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09339_ _10172_/A1 _09343_/B _08851_/A vssd1 vssd1 vccd1 vccd1 _09339_/X sky130_fd_sc_hd__a21o_1
XFILLER_55_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11301_ _11332_/CLK _11301_/D vssd1 vssd1 vccd1 vccd1 _11301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11232_ _11651_/CLK _11232_/D vssd1 vssd1 vccd1 vccd1 _11232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11163_ _11683_/CLK _11163_/D vssd1 vssd1 vccd1 vccd1 _11163_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11762_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10114_ _10114_/A0 _11761_/Q _10118_/S vssd1 vssd1 vccd1 vccd1 _11761_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11094_ _11312_/CLK _11094_/D vssd1 vssd1 vccd1 vccd1 _11094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10045_ _11714_/Q _07070_/A _10051_/S vssd1 vssd1 vccd1 vccd1 _10046_/B sky130_fd_sc_hd__mux2_1
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10947_ _11023_/CLK _10947_/D vssd1 vssd1 vccd1 vccd1 _10947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10878_ _10929_/CLK _10878_/D vssd1 vssd1 vccd1 vccd1 _10878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_2 _05259_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout509 fanout510/X vssd1 vssd1 vccd1 vccd1 _09048_/C1 sky130_fd_sc_hd__buf_4
XFILLER_141_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _08956_/B _09668_/C vssd1 vssd1 vccd1 vccd1 _06971_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08710_ _08810_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _11209_/D sky130_fd_sc_hd__or2_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05922_ _05922_/A _05922_/B _05922_/C vssd1 vssd1 vccd1 vccd1 _05922_/X sky130_fd_sc_hd__and3_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09690_ _05396_/S _09682_/B _09682_/Y _11637_/Q _09689_/X vssd1 vssd1 vccd1 vccd1
+ _09691_/B sky130_fd_sc_hd__o221a_1
XFILLER_94_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08641_ _11175_/Q _08645_/S _07086_/Y _07005_/A vssd1 vssd1 vccd1 vccd1 _11175_/D
+ sky130_fd_sc_hd__o22a_1
X_05853_ _10397_/Q _06804_/B _06805_/B1 _10533_/Q _05850_/X vssd1 vssd1 vccd1 vccd1
+ _05853_/X sky130_fd_sc_hd__o221a_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08572_ _11141_/Q _08834_/A0 _08577_/S vssd1 vssd1 vccd1 vccd1 _08573_/B sky130_fd_sc_hd__mux2_1
X_05784_ _10697_/Q _06807_/A2 _05780_/X _05783_/X vssd1 vssd1 vccd1 vccd1 _05784_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_81_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07523_ _08423_/A1 _10546_/Q _07535_/S vssd1 vssd1 vccd1 vccd1 _07524_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07454_ _07455_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07752_/B sky130_fd_sc_hd__nor2_4
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06405_ _07690_/A _06404_/X _06403_/X _07082_/A vssd1 vssd1 vccd1 vccd1 _06405_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_50_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07385_ _10468_/Q _10128_/A0 _07393_/S vssd1 vssd1 vccd1 vccd1 _07386_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09124_ _09124_/A1 _09110_/X _09123_/X _09279_/C1 vssd1 vssd1 vccd1 vccd1 _11408_/D
+ sky130_fd_sc_hd__o211a_1
X_06336_ _11215_/Q _06126_/B _06332_/X _06335_/X vssd1 vssd1 vccd1 vccd1 _06336_/X
+ sky130_fd_sc_hd__o211a_1
X_09055_ _11377_/Q _09055_/B vssd1 vssd1 vccd1 vccd1 _09055_/X sky130_fd_sc_hd__or2_1
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06267_ _10872_/Q _06318_/A2 _06453_/B1 _10990_/Q vssd1 vssd1 vccd1 vccd1 _06267_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05218_ _11056_/Q _11055_/Q _11595_/Q vssd1 vssd1 vccd1 vccd1 _05223_/B sky130_fd_sc_hd__mux2_1
XFILLER_85_1311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08006_ _10190_/A0 _08011_/S _08005_/X _08351_/C1 vssd1 vssd1 vccd1 vccd1 _10827_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06198_ _10284_/Q _06106_/B _06197_/X _06997_/A vssd1 vssd1 vccd1 vccd1 _06198_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05149_ _10938_/Q _10937_/Q _05429_/S vssd1 vssd1 vccd1 vccd1 _05151_/C sky130_fd_sc_hd__mux2_1
XFILLER_131_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09957_ _09957_/A _09957_/B _09957_/C _09957_/D vssd1 vssd1 vccd1 vccd1 _09958_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08908_ _11313_/Q _08946_/B vssd1 vssd1 vccd1 vccd1 _08908_/X sky130_fd_sc_hd__or2_1
XFILLER_58_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09888_ _09908_/A _09888_/B _09888_/C vssd1 vssd1 vccd1 vccd1 _09889_/A sky130_fd_sc_hd__or3_2
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _08839_/A _08839_/B vssd1 vssd1 vccd1 vccd1 _11277_/D sky130_fd_sc_hd__or2_1
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_tms1x00_1101 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1101/HI io_oeb[31] sky130_fd_sc_hd__conb_1
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_tms1x00_1112 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1112/HI io_out[4] sky130_fd_sc_hd__conb_1
XFILLER_131_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1123 vssd1 vssd1 vccd1 vccd1 io_oeb[0] wrapped_tms1x00_1123/LO sky130_fd_sc_hd__conb_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10801_ _11698_/CLK _10801_/D vssd1 vssd1 vccd1 vccd1 _10801_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _11781_/CLK _11781_/D vssd1 vssd1 vccd1 vccd1 _11781_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10732_ _11706_/CLK _10732_/D vssd1 vssd1 vccd1 vccd1 _10732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10663_ _11458_/CLK _10663_/D vssd1 vssd1 vccd1 vccd1 _10663_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10594_ _11280_/CLK _10594_/D vssd1 vssd1 vccd1 vccd1 _10594_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_154_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11215_ _11220_/CLK _11215_/D vssd1 vssd1 vccd1 vccd1 _11215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11146_ _11151_/CLK _11146_/D vssd1 vssd1 vccd1 vccd1 _11146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11077_ _11768_/CLK _11077_/D vssd1 vssd1 vccd1 vccd1 _11077_/Q sky130_fd_sc_hd__dfxtp_1
X_10028_ _10028_/A _10028_/B vssd1 vssd1 vccd1 vccd1 _10085_/S sky130_fd_sc_hd__nand2_8
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07170_ _08846_/A0 _10346_/Q _09243_/C vssd1 vssd1 vccd1 vccd1 _07171_/B sky130_fd_sc_hd__mux2_1
XFILLER_121_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06121_ _11224_/Q _07190_/A _06373_/B1 _10813_/Q vssd1 vssd1 vccd1 vccd1 _06125_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06052_ _11037_/Q _08383_/A _09154_/A _11193_/Q _06051_/X vssd1 vssd1 vccd1 vccd1
+ _06052_/X sky130_fd_sc_hd__o221a_1
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout306 _07751_/A2 vssd1 vssd1 vccd1 vccd1 _07761_/A2 sky130_fd_sc_hd__clkbuf_8
X_09811_ _09811_/A _09811_/B _09811_/C _09811_/D vssd1 vssd1 vccd1 vccd1 _09811_/X
+ sky130_fd_sc_hd__or4_1
Xfanout317 _07977_/S vssd1 vssd1 vccd1 vccd1 _07991_/S sky130_fd_sc_hd__buf_8
XFILLER_115_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout328 _07425_/S vssd1 vssd1 vccd1 vccd1 _07437_/S sky130_fd_sc_hd__buf_8
XFILLER_115_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout339 _09426_/S vssd1 vssd1 vccd1 vccd1 _09704_/B sky130_fd_sc_hd__buf_8
XFILLER_98_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09742_ _10504_/Q _09568_/A _09874_/A2 _10496_/Q _09741_/X vssd1 vssd1 vccd1 vccd1
+ _09749_/A sky130_fd_sc_hd__a221o_1
X_06954_ _06944_/Y _09538_/D _11606_/Q _09538_/C vssd1 vssd1 vccd1 vccd1 _06954_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05905_ _10258_/Q _06976_/A _06351_/A2 _10205_/Q _05904_/X vssd1 vssd1 vccd1 vccd1
+ _05905_/X sky130_fd_sc_hd__o221a_1
XFILLER_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09673_ _11629_/Q _09673_/B vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__nand2_8
X_06885_ _09395_/A0 _07048_/A _08970_/S _06884_/Y _10217_/Q vssd1 vssd1 vccd1 vccd1
+ _10217_/D sky130_fd_sc_hd__a32o_1
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _08941_/A _08624_/B vssd1 vssd1 vccd1 vccd1 _11166_/D sky130_fd_sc_hd__or2_1
X_05836_ _11667_/Q _09965_/A _09314_/A _11509_/Q _05835_/X vssd1 vssd1 vccd1 vccd1
+ _05836_/X sky130_fd_sc_hd__o221a_1
XFILLER_43_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05767_ _11756_/Q _10108_/A _05763_/X _05766_/X vssd1 vssd1 vccd1 vccd1 _05767_/X
+ sky130_fd_sc_hd__o211a_4
X_08555_ _11131_/Q _08558_/S _07357_/S _07314_/B vssd1 vssd1 vccd1 vccd1 _11131_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07506_ _07790_/A _07506_/B vssd1 vssd1 vccd1 vccd1 _10537_/D sky130_fd_sc_hd__or2_1
XFILLER_23_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05698_ _11116_/Q _05615_/Y _05621_/Y _11115_/Q _05697_/X vssd1 vssd1 vccd1 vccd1
+ _05703_/A sky130_fd_sc_hd__a221o_1
X_08486_ _10115_/A0 _08497_/S _08485_/X _09022_/C1 vssd1 vssd1 vccd1 vccd1 _11093_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07437_ _07036_/A _10495_/Q _07437_/S vssd1 vssd1 vccd1 vccd1 _07438_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07368_ _10456_/Q _08326_/B2 _07373_/S vssd1 vssd1 vccd1 vccd1 _10456_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09107_ _11401_/Q _09243_/B _07591_/S _09192_/A vssd1 vssd1 vccd1 vccd1 _09107_/X
+ sky130_fd_sc_hd__a31o_1
X_06319_ _10587_/Q _06539_/A2 _06539_/B1 _10838_/Q _06624_/C1 vssd1 vssd1 vccd1 vccd1
+ _06319_/X sky130_fd_sc_hd__o221a_1
XFILLER_136_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07299_ _09325_/A _08471_/B _10136_/C vssd1 vssd1 vccd1 vccd1 _08762_/B sky130_fd_sc_hd__and3_4
X_09038_ _09038_/A _09271_/B _09038_/C vssd1 vssd1 vccd1 vccd1 _09038_/X sky130_fd_sc_hd__or3_4
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11000_ _11675_/CLK _11000_/D vssd1 vssd1 vccd1 vccd1 _11000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout840 _06861_/B vssd1 vssd1 vccd1 vccd1 _07853_/A sky130_fd_sc_hd__buf_6
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout851 fanout861/X vssd1 vssd1 vccd1 vccd1 _06642_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_120_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout862 _06871_/A2 vssd1 vssd1 vccd1 vccd1 _06860_/A2 sky130_fd_sc_hd__buf_6
Xfanout873 _05741_/Y vssd1 vssd1 vccd1 vccd1 _06719_/A2 sky130_fd_sc_hd__buf_8
Xfanout884 _06227_/A2 vssd1 vssd1 vccd1 vccd1 _09998_/A sky130_fd_sc_hd__buf_6
XFILLER_93_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout895 fanout901/X vssd1 vssd1 vccd1 vccd1 _06539_/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_200 _10021_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11765_/CLK _11764_/D vssd1 vssd1 vccd1 vccd1 _11764_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10785_/CLK _10715_/D vssd1 vssd1 vccd1 vccd1 _10715_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11695_ _11765_/CLK _11695_/D vssd1 vssd1 vccd1 vccd1 _11695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10646_ _11270_/CLK _10646_/D vssd1 vssd1 vccd1 vccd1 _10646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10577_ _10808_/CLK _10577_/D vssd1 vssd1 vccd1 vccd1 _10577_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_51_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11186_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11129_ _11268_/CLK _11129_/D vssd1 vssd1 vccd1 vccd1 _11129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06670_ _10487_/Q _06872_/A2 _06667_/X _06669_/X _06670_/D1 vssd1 vssd1 vccd1 vccd1
+ _06670_/X sky130_fd_sc_hd__o2111a_1
XFILLER_149_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05621_ _05621_/A _05621_/B vssd1 vssd1 vccd1 vccd1 _05621_/Y sky130_fd_sc_hd__nor2_8
XFILLER_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05552_ _05618_/A1 _11425_/Q _11422_/Q _05606_/B2 _05550_/X vssd1 vssd1 vccd1 vccd1
+ _05555_/A sky130_fd_sc_hd__a221o_4
X_08340_ _11013_/Q _08362_/B vssd1 vssd1 vccd1 vccd1 _08340_/X sky130_fd_sc_hd__or2_1
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08271_ _08846_/A0 _08272_/S _08270_/X _08791_/C1 vssd1 vssd1 vccd1 vccd1 _10967_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05483_ _10228_/Q input70/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05483_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07222_ _07222_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _07222_/Y sky130_fd_sc_hd__nor2_4
XFILLER_118_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07153_ _07153_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _09240_/S sky130_fd_sc_hd__or2_4
XFILLER_34_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06104_ _06189_/A1 _06098_/X _06103_/X _08243_/A _06093_/X vssd1 vssd1 vccd1 vccd1
+ _06104_/X sky130_fd_sc_hd__o311a_2
X_07084_ _07689_/A _07690_/B vssd1 vssd1 vccd1 vccd1 _10108_/C sky130_fd_sc_hd__nand2_1
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06035_ _11363_/Q _09016_/A _08994_/A _11353_/Q _06349_/C1 vssd1 vssd1 vccd1 vccd1
+ _06035_/X sky130_fd_sc_hd__o221a_1
XFILLER_82_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07986_ _10818_/Q _10132_/A0 _07991_/S vssd1 vssd1 vccd1 vccd1 _07987_/B sky130_fd_sc_hd__mux2_1
X_09725_ _10342_/Q _09873_/A2 _09873_/B1 _10347_/Q vssd1 vssd1 vccd1 vccd1 _09725_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06937_ _10213_/Q _06937_/B vssd1 vssd1 vccd1 vccd1 _08950_/B sky130_fd_sc_hd__nand2_8
XFILLER_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09656_ _10337_/Q _09572_/A _09950_/B1 _10318_/Q _09655_/X vssd1 vssd1 vccd1 vccd1
+ _09659_/C sky130_fd_sc_hd__a221o_1
XFILLER_103_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06868_ _06883_/B _06868_/B vssd1 vssd1 vccd1 vccd1 _10250_/D sky130_fd_sc_hd__and2_1
XFILLER_43_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _09285_/A1 _11158_/Q _08623_/S vssd1 vssd1 vccd1 vccd1 _08608_/B sky130_fd_sc_hd__mux2_1
X_05819_ _05819_/A _05819_/B vssd1 vssd1 vccd1 vccd1 _05819_/Y sky130_fd_sc_hd__nor2_8
XFILLER_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _10273_/Q _09565_/A _09570_/B _10274_/Q vssd1 vssd1 vccd1 vccd1 _09587_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ _10696_/Q _06799_/A2 _06870_/B1 _10520_/Q vssd1 vssd1 vccd1 vccd1 _06799_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08684_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _11118_/D sky130_fd_sc_hd__or2_1
XFILLER_24_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08469_ _08469_/A _08469_/B _10180_/C _10119_/B vssd1 vssd1 vccd1 vccd1 _08469_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10500_ _11470_/CLK _10500_/D vssd1 vssd1 vccd1 vccd1 _10500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11480_ _11685_/CLK _11480_/D vssd1 vssd1 vccd1 vccd1 _11480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10431_ _11284_/CLK _10431_/D vssd1 vssd1 vccd1 vccd1 _10431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10362_ _11722_/CLK _10362_/D vssd1 vssd1 vccd1 vccd1 _10362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10293_ _11719_/CLK _10293_/D vssd1 vssd1 vccd1 vccd1 _10293_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout670 _06942_/A vssd1 vssd1 vccd1 vccd1 _05471_/A sky130_fd_sc_hd__buf_8
XFILLER_59_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout681 _05432_/S vssd1 vssd1 vccd1 vccd1 _05377_/S sky130_fd_sc_hd__buf_8
Xfanout692 _11596_/Q vssd1 vssd1 vccd1 vccd1 _05372_/S sky130_fd_sc_hd__buf_12
XFILLER_98_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11809_/CLK _11747_/D vssd1 vssd1 vccd1 vccd1 _11747_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _11684_/CLK _11678_/D vssd1 vssd1 vccd1 vccd1 _11678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10629_ _11703_/CLK _10629_/D vssd1 vssd1 vccd1 vccd1 _10629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07840_ _07143_/A _07819_/Y _07961_/S _10735_/Q vssd1 vssd1 vccd1 vccd1 _10735_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07771_ _07335_/B _07204_/B _07771_/B1 _10691_/Q _07309_/A vssd1 vssd1 vccd1 vccd1
+ _10691_/D sky130_fd_sc_hd__a221o_1
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09510_ _09492_/B _09502_/B _09508_/Y _09509_/X _09529_/A vssd1 vssd1 vccd1 vccd1
+ _11613_/D sky130_fd_sc_hd__o311a_1
X_06722_ _06855_/B _06715_/Y _06720_/Y _06721_/Y vssd1 vssd1 vccd1 vccd1 _06722_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_83_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _09441_/A _09441_/B vssd1 vssd1 vccd1 vccd1 _09441_/Y sky130_fd_sc_hd__nor2_2
X_06653_ _10358_/Q _08649_/A _06651_/X _06652_/X vssd1 vssd1 vccd1 vccd1 _06653_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05604_ _05628_/A2 _11545_/Q _11542_/Q _05628_/B1 vssd1 vssd1 vccd1 vccd1 _05604_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09372_ _10172_/A1 _09376_/B _10178_/B1 vssd1 vssd1 vccd1 vccd1 _09372_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06584_ _11031_/Q _09016_/A _06580_/X _06583_/X vssd1 vssd1 vccd1 vccd1 _06584_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08323_ _08323_/A _08325_/B vssd1 vssd1 vccd1 vccd1 _08323_/Y sky130_fd_sc_hd__nand2_1
X_05535_ _05631_/A2 _11527_/Q _11523_/Q _05631_/B1 _05533_/X vssd1 vssd1 vccd1 vccd1
+ _05535_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05466_ _05466_/A _05466_/B _05466_/C _05466_/D vssd1 vssd1 vccd1 vccd1 _05470_/A
+ sky130_fd_sc_hd__or4_1
X_08254_ _09141_/A1 _10959_/Q _08272_/S vssd1 vssd1 vccd1 vccd1 _08255_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07205_ _07205_/A _07205_/B vssd1 vssd1 vccd1 vccd1 _07205_/Y sky130_fd_sc_hd__nand2_2
XFILLER_118_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05397_ _11218_/Q _11217_/Q _05397_/S vssd1 vssd1 vccd1 vccd1 _05400_/B sky130_fd_sc_hd__mux2_1
X_08185_ _08810_/A _08185_/B vssd1 vssd1 vccd1 vccd1 _10926_/D sky130_fd_sc_hd__or2_1
XFILLER_152_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07136_ _10329_/Q _07145_/B vssd1 vssd1 vccd1 vccd1 _07136_/X sky130_fd_sc_hd__or2_1
XFILLER_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07067_ _10292_/Q _07078_/B _07496_/S _07241_/B vssd1 vssd1 vccd1 vccd1 _10292_/D
+ sky130_fd_sc_hd__o22a_1
X_06018_ _11522_/Q _09326_/A _06363_/A2 _11482_/Q vssd1 vssd1 vccd1 vccd1 _06018_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_88_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07969_ _10807_/Q _07441_/A _07901_/B _07968_/X vssd1 vssd1 vccd1 vccd1 _10807_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_114_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09708_ _10396_/Q _09874_/A2 _09873_/B1 _10405_/Q _09707_/X vssd1 vssd1 vccd1 vccd1
+ _09713_/B sky130_fd_sc_hd__a221o_1
X_10980_ _10981_/CLK _10980_/D vssd1 vssd1 vccd1 vccd1 _10980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09639_ _09600_/B _09561_/B _09637_/X _09638_/Y _09827_/A vssd1 vssd1 vccd1 vccd1
+ _09640_/C sky130_fd_sc_hd__o221a_1
XFILLER_83_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11601_ _11601_/CLK _11601_/D vssd1 vssd1 vccd1 vccd1 _11601_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11532_ _11762_/CLK _11532_/D vssd1 vssd1 vccd1 vccd1 _11532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11463_ _11473_/CLK _11463_/D vssd1 vssd1 vccd1 vccd1 _11463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10414_ _11458_/CLK _10414_/D vssd1 vssd1 vccd1 vccd1 _10414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11394_ _11410_/CLK _11394_/D vssd1 vssd1 vccd1 vccd1 _11394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10345_ _10765_/CLK _10345_/D vssd1 vssd1 vccd1 vccd1 _10345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10276_ _11710_/CLK _10276_/D vssd1 vssd1 vccd1 vccd1 _10276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05320_ _10885_/Q _10884_/Q _05397_/S vssd1 vssd1 vccd1 vccd1 _05323_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05251_ _10980_/Q _10979_/Q _05382_/S vssd1 vssd1 vccd1 vccd1 _05253_/C sky130_fd_sc_hd__mux2_1
XFILLER_70_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05182_ _10592_/Q _10835_/Q _06939_/A vssd1 vssd1 vccd1 vccd1 _05184_/C sky130_fd_sc_hd__mux2_1
XFILLER_31_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09990_ _10172_/A1 _09994_/B _08618_/A vssd1 vssd1 vccd1 vccd1 _09990_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08941_ _08941_/A _08941_/B vssd1 vssd1 vccd1 vccd1 _11329_/D sky130_fd_sc_hd__or2_1
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08872_ _09172_/A1 _11293_/Q _08890_/S vssd1 vssd1 vccd1 vccd1 _08873_/B sky130_fd_sc_hd__mux2_1
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07823_ _07007_/A _07839_/A2 _07821_/A _10718_/Q vssd1 vssd1 vccd1 vccd1 _10718_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07754_ _10678_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07754_/X sky130_fd_sc_hd__or2_1
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06705_ _11445_/Q _07777_/A _06875_/A2 _10781_/Q vssd1 vssd1 vccd1 vccd1 _06705_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07685_ _10641_/Q _07673_/Y _07676_/X _09232_/B2 vssd1 vssd1 vccd1 vccd1 _10641_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09424_ _11640_/Q _11583_/Q _09704_/B vssd1 vssd1 vccd1 vccd1 _11583_/D sky130_fd_sc_hd__mux2_1
X_06636_ _11080_/Q _06636_/A2 _05865_/B _11781_/Q _06635_/X vssd1 vssd1 vccd1 vccd1
+ _06636_/X sky130_fd_sc_hd__o221a_1
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09355_ _10080_/A0 _11535_/Q _09357_/S vssd1 vssd1 vccd1 vccd1 _11535_/D sky130_fd_sc_hd__mux2_1
X_06567_ _11708_/Q _08560_/A _06565_/X _06566_/X vssd1 vssd1 vccd1 vccd1 _06567_/X
+ sky130_fd_sc_hd__a211o_1
X_08306_ _10986_/Q _08302_/Y _08303_/Y _08441_/B2 vssd1 vssd1 vccd1 vccd1 _10986_/D
+ sky130_fd_sc_hd__o22a_1
X_05518_ _05518_/A _05518_/B vssd1 vssd1 vccd1 vccd1 _05518_/Y sky130_fd_sc_hd__nor2_8
X_09286_ _10023_/A0 _09288_/B _09290_/B1 vssd1 vssd1 vccd1 vccd1 _09286_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06498_ _10945_/Q _06630_/A2 _06630_/B1 _11021_/Q vssd1 vssd1 vccd1 vccd1 _06498_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08237_ _10952_/Q _08324_/B vssd1 vssd1 vccd1 vccd1 _08237_/X sky130_fd_sc_hd__or2_1
X_05449_ _05449_/A _05449_/B _05449_/C _05449_/D vssd1 vssd1 vccd1 vccd1 _05452_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_14_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08168_ _07002_/A _10910_/Q _08182_/S vssd1 vssd1 vccd1 vccd1 _10910_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_108_wb_clk_i clkbuf_4_10__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11458_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07119_ _10316_/Q _07145_/B _07188_/S _07095_/B vssd1 vssd1 vccd1 vccd1 _10316_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_84_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08099_ _08092_/X _08354_/S _08098_/X _08427_/A vssd1 vssd1 vccd1 vccd1 _10873_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10130_ _07059_/A _11776_/Q _10134_/S vssd1 vssd1 vccd1 vccd1 _11776_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10061_ _10061_/A _10108_/B _10119_/C vssd1 vssd1 vccd1 vccd1 _10071_/S sky130_fd_sc_hd__or3_4
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10963_ _11243_/CLK _10963_/D vssd1 vssd1 vccd1 vccd1 _10963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10894_ _11632_/CLK _10894_/D vssd1 vssd1 vccd1 vccd1 _10894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11515_ _11735_/CLK _11515_/D vssd1 vssd1 vccd1 vccd1 _11515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ _11450_/CLK _11446_/D vssd1 vssd1 vccd1 vccd1 _11446_/Q sky130_fd_sc_hd__dfxtp_1
X_11377_ _11497_/CLK _11377_/D vssd1 vssd1 vccd1 vccd1 _11377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _10725_/CLK _10328_/D vssd1 vssd1 vccd1 vccd1 _10328_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10259_ _11755_/CLK _10259_/D vssd1 vssd1 vccd1 vccd1 _10259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07470_ _07476_/A _07470_/B vssd1 vssd1 vccd1 vccd1 _10512_/D sky130_fd_sc_hd__or2_1
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06421_ _10919_/Q _06591_/A2 _06126_/B _10744_/Q vssd1 vssd1 vccd1 vccd1 _06421_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_50_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09140_ _09985_/A1 _09132_/X _09139_/X _10175_/C1 vssd1 vssd1 vccd1 vccd1 _11415_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06352_ _11811_/Q _10180_/A _06348_/X _06351_/X vssd1 vssd1 vccd1 vccd1 _06353_/C
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11584_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05303_ _11020_/Q _11019_/Q _05413_/S vssd1 vssd1 vccd1 vccd1 _05307_/A sky130_fd_sc_hd__mux2_1
X_06283_ _11810_/Q _10180_/A _08097_/A _10201_/Q vssd1 vssd1 vccd1 vccd1 _06283_/X
+ sky130_fd_sc_hd__o22a_1
X_09071_ _09283_/A1 _09077_/B _08783_/A vssd1 vssd1 vccd1 vccd1 _09071_/X sky130_fd_sc_hd__a21o_1
X_08022_ _09364_/A1 _08035_/S _08021_/X _07011_/B vssd1 vssd1 vccd1 vccd1 _10835_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05234_ _05471_/A _10953_/Q vssd1 vssd1 vccd1 vccd1 _05234_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05165_ _11074_/Q _11073_/Q _05393_/S vssd1 vssd1 vccd1 vccd1 _05167_/C sky130_fd_sc_hd__mux2_1
XFILLER_116_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09973_ _10080_/A0 _11673_/Q _09975_/S vssd1 vssd1 vccd1 vccd1 _11673_/D sky130_fd_sc_hd__mux2_1
X_05096_ _11872_/A vssd1 vssd1 vccd1 vccd1 _08243_/B sky130_fd_sc_hd__inv_8
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08924_ _11321_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08924_/X sky130_fd_sc_hd__or2_1
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08855_ _08855_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08855_/X sky130_fd_sc_hd__or2_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07806_ _07922_/A _07806_/B vssd1 vssd1 vccd1 vccd1 _10710_/D sky130_fd_sc_hd__or2_1
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08786_ _08876_/A0 _11249_/Q _08802_/S vssd1 vssd1 vccd1 vccd1 _08787_/B sky130_fd_sc_hd__mux2_1
X_05998_ _11210_/Q _06126_/B _05996_/X _05997_/X vssd1 vssd1 vccd1 vccd1 _05998_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _07025_/A _07761_/A2 _07736_/X _09201_/A1 vssd1 vssd1 vccd1 vccd1 _10669_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07668_ _10629_/Q _07665_/S _07233_/S _07187_/B vssd1 vssd1 vccd1 vccd1 _10629_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09407_ _09407_/A _09407_/B vssd1 vssd1 vccd1 vccd1 _09414_/S sky130_fd_sc_hd__nand2_8
XFILLER_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06619_ _06619_/A1 _06590_/X _06601_/X _06618_/X vssd1 vssd1 vccd1 vccd1 _06619_/X
+ sky130_fd_sc_hd__a31o_1
X_07599_ _07599_/A _08852_/B vssd1 vssd1 vccd1 vccd1 _07599_/Y sky130_fd_sc_hd__nor2_2
XFILLER_71_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09338_ _11523_/Q _09326_/X _09337_/X vssd1 vssd1 vccd1 vccd1 _11523_/D sky130_fd_sc_hd__a21o_1
XFILLER_90_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09269_ _11487_/Q _09249_/X _09268_/X vssd1 vssd1 vccd1 vccd1 _11487_/D sky130_fd_sc_hd__a21o_1
X_11300_ _11325_/CLK _11300_/D vssd1 vssd1 vccd1 vccd1 _11300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11231_ _11652_/CLK _11231_/D vssd1 vssd1 vccd1 vccd1 _11231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11162_ _11332_/CLK _11162_/D vssd1 vssd1 vccd1 vccd1 _11162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10113_ _10113_/A0 _11760_/Q _10118_/S vssd1 vssd1 vccd1 vccd1 _11760_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11093_ _11811_/CLK _11093_/D vssd1 vssd1 vccd1 vccd1 _11093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10044_ _11713_/Q _10028_/B _10085_/S _07243_/B vssd1 vssd1 vccd1 vccd1 _11713_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_76_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11393_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10946_ _11733_/CLK _10946_/D vssd1 vssd1 vccd1 vccd1 _10946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10877_ _10929_/CLK _10877_/D vssd1 vssd1 vccd1 vccd1 _10877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 _05259_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11429_ _11801_/CLK _11429_/D vssd1 vssd1 vccd1 vccd1 _11429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ input9/X _09668_/C vssd1 vssd1 vccd1 vccd1 _06970_/X sky130_fd_sc_hd__and2_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05921_ _11105_/Q _09082_/A _06697_/B1 _11241_/Q vssd1 vssd1 vccd1 vccd1 _05922_/C
+ sky130_fd_sc_hd__o22a_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1070 _10142_/A1 vssd1 vssd1 vccd1 vccd1 _10015_/A0 sky130_fd_sc_hd__buf_6
XFILLER_55_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08640_ _07232_/B _08637_/C _08639_/X vssd1 vssd1 vccd1 vccd1 _11174_/D sky130_fd_sc_hd__a21o_1
X_05852_ _10698_/Q _06807_/A2 _07540_/A _10555_/Q _05849_/X vssd1 vssd1 vccd1 vccd1
+ _05852_/X sky130_fd_sc_hd__o221a_2
XFILLER_94_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08571_ _11140_/Q _08577_/S _08563_/Y _07098_/B vssd1 vssd1 vccd1 vccd1 _11140_/D
+ sky130_fd_sc_hd__o22a_1
X_05783_ _11451_/Q _06194_/A2 _05782_/X _06808_/C1 vssd1 vssd1 vccd1 vccd1 _05783_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07522_ _07926_/A _07522_/B vssd1 vssd1 vccd1 vccd1 _10545_/D sky130_fd_sc_hd__or2_1
XFILLER_74_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07453_ _10504_/Q _07441_/Y _07443_/Y _07040_/X vssd1 vssd1 vccd1 vccd1 _10504_/D
+ sky130_fd_sc_hd__a22o_1
X_06404_ _06388_/X _06389_/X _06392_/X _06387_/X vssd1 vssd1 vccd1 vccd1 _06404_/X
+ sky130_fd_sc_hd__a31o_1
X_07384_ _10467_/Q _07380_/S _07655_/S _07232_/B vssd1 vssd1 vccd1 vccd1 _10467_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09123_ _11408_/Q _09127_/B vssd1 vssd1 vccd1 vccd1 _09123_/X sky130_fd_sc_hd__or2_1
XFILLER_109_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06335_ _11263_/Q _06635_/B1 _06333_/X _06334_/X vssd1 vssd1 vccd1 vccd1 _06335_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09054_ _11376_/Q _09038_/X _09053_/X vssd1 vssd1 vccd1 vccd1 _11376_/D sky130_fd_sc_hd__a21o_1
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06266_ _10864_/Q _06540_/A2 _06262_/X _06265_/X vssd1 vssd1 vccd1 vccd1 _06266_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08005_ _10827_/Q _08091_/C vssd1 vssd1 vccd1 vccd1 _08005_/X sky130_fd_sc_hd__or2_1
X_05217_ _10858_/Q _10857_/Q _09680_/C vssd1 vssd1 vccd1 vccd1 _05223_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06197_ _10316_/Q _06856_/A2 _06710_/B _10720_/Q _06196_/X vssd1 vssd1 vccd1 vccd1
+ _06197_/X sky130_fd_sc_hd__o221a_1
XFILLER_85_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05148_ _11312_/Q _11311_/Q _05426_/S vssd1 vssd1 vccd1 vccd1 _05151_/B sky130_fd_sc_hd__mux2_1
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05079_ _05079_/A vssd1 vssd1 vccd1 vccd1 _05079_/Y sky130_fd_sc_hd__inv_2
X_09956_ _10696_/Q _09571_/A _09573_/D _10687_/Q vssd1 vssd1 vccd1 vccd1 _09957_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08907_ _08907_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08907_/X sky130_fd_sc_hd__or2_2
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09887_/A _09887_/B _09887_/C _09887_/D vssd1 vssd1 vccd1 vccd1 _09888_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _08838_/A0 _11277_/Q _08838_/S vssd1 vssd1 vccd1 vccd1 _08839_/B sky130_fd_sc_hd__mux2_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1102 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1102/HI io_oeb[32] sky130_fd_sc_hd__conb_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1113 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1113/HI io_out[5] sky130_fd_sc_hd__conb_1
XFILLER_79_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1124 vssd1 vssd1 vccd1 vccd1 io_oeb[1] wrapped_tms1x00_1124/LO sky130_fd_sc_hd__conb_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _08869_/A _08769_/B vssd1 vssd1 vccd1 vccd1 _11240_/D sky130_fd_sc_hd__or2_1
XFILLER_22_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _11743_/CLK _10800_/D vssd1 vssd1 vccd1 vccd1 _10800_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11780_/CLK _11780_/D vssd1 vssd1 vccd1 vccd1 _11780_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10731_ _11719_/CLK _10731_/D vssd1 vssd1 vccd1 vccd1 _10731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10662_ _10785_/CLK _10662_/D vssd1 vssd1 vccd1 vccd1 _10662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_123_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11713_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10593_ _11243_/CLK _10593_/D vssd1 vssd1 vccd1 vccd1 _10593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ _11770_/CLK _11214_/D vssd1 vssd1 vccd1 vccd1 _11214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11145_ _11151_/CLK _11145_/D vssd1 vssd1 vccd1 vccd1 _11145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11076_ _11268_/CLK _11076_/D vssd1 vssd1 vccd1 vccd1 _11076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10027_ _10039_/A _10051_/S vssd1 vssd1 vccd1 vccd1 _10027_/Y sky130_fd_sc_hd__nor2_2
XFILLER_97_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10929_ _10929_/CLK _10929_/D vssd1 vssd1 vccd1 vccd1 _10929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06120_ _11194_/Q _06736_/A2 _06221_/A2 _11157_/Q _06119_/X vssd1 vssd1 vccd1 vccd1
+ _06120_/X sky130_fd_sc_hd__o221a_4
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06051_ _10959_/Q _06363_/A2 _09132_/A _11289_/Q vssd1 vssd1 vccd1 vccd1 _06051_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09810_ _10280_/Q _09566_/A _09568_/D _10281_/Q _09805_/X vssd1 vssd1 vccd1 vccd1
+ _09811_/D sky130_fd_sc_hd__a221o_1
Xfanout307 _07455_/X vssd1 vssd1 vccd1 vccd1 _07751_/A2 sky130_fd_sc_hd__buf_6
Xfanout318 _07353_/B vssd1 vssd1 vccd1 vccd1 _08558_/S sky130_fd_sc_hd__buf_6
XFILLER_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout329 _07190_/X vssd1 vssd1 vccd1 vccd1 _07425_/S sky130_fd_sc_hd__buf_8
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09741_ _10542_/Q _09873_/B1 _09875_/B1 _10533_/Q vssd1 vssd1 vccd1 vccd1 _09741_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_101_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06953_ _09539_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09538_/D sky130_fd_sc_hd__nor2_2
XFILLER_80_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05904_ _11361_/Q _09016_/A _08472_/A _11351_/Q _07689_/B vssd1 vssd1 vccd1 vccd1
+ _05904_/X sky130_fd_sc_hd__o221a_1
XFILLER_100_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09672_ _11629_/Q _09672_/B vssd1 vssd1 vccd1 vccd1 _09672_/Y sky130_fd_sc_hd__nor2_2
XFILLER_80_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06884_ input74/X _08970_/S vssd1 vssd1 vccd1 vccd1 _06884_/Y sky130_fd_sc_hd__nor2_4
XFILLER_95_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08623_ _08937_/A1 _11166_/Q _08623_/S vssd1 vssd1 vccd1 vccd1 _08624_/B sky130_fd_sc_hd__mux2_1
X_05835_ _11724_/Q _08200_/A _08097_/A _11529_/Q vssd1 vssd1 vccd1 vccd1 _05835_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08554_ _11130_/Q _08558_/S _07355_/S _08811_/B2 vssd1 vssd1 vccd1 vccd1 _11130_/D
+ sky130_fd_sc_hd__o22a_1
X_05766_ _11508_/Q _09314_/A _05764_/X _05765_/X vssd1 vssd1 vccd1 vccd1 _05766_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07505_ _10023_/A0 _10537_/Q _07513_/S vssd1 vssd1 vccd1 vccd1 _07506_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08485_ _11093_/Q _08503_/B vssd1 vssd1 vccd1 vccd1 _08485_/X sky130_fd_sc_hd__or2_1
X_05697_ _11120_/Q _05543_/Y _05603_/Y _11107_/Q vssd1 vssd1 vccd1 vccd1 _05697_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07436_ _10058_/A _07436_/B vssd1 vssd1 vccd1 vccd1 _10494_/D sky130_fd_sc_hd__or2_1
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07367_ _10455_/Q _07088_/X _07373_/S vssd1 vssd1 vccd1 vccd1 _10455_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09106_ _07040_/B _07539_/Y _09105_/X vssd1 vssd1 vccd1 vccd1 _11400_/D sky130_fd_sc_hd__a21o_1
X_06318_ _10423_/Q _06318_/A2 _06453_/B1 _10641_/Q vssd1 vssd1 vccd1 vccd1 _06318_/X
+ sky130_fd_sc_hd__o22a_1
X_07298_ _07689_/A _07298_/B vssd1 vssd1 vccd1 vccd1 _07298_/X sky130_fd_sc_hd__or2_1
XFILLER_136_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09037_ _09037_/A _10136_/B _09037_/C vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__and3_4
X_06249_ _11292_/Q _06739_/A2 _06718_/C1 _06248_/X vssd1 vssd1 vccd1 vccd1 _06249_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout830 _06161_/A2 vssd1 vssd1 vccd1 vccd1 _10108_/A sky130_fd_sc_hd__buf_6
Xfanout841 fanout846/X vssd1 vssd1 vccd1 vccd1 _06861_/B sky130_fd_sc_hd__buf_6
Xfanout852 fanout861/X vssd1 vssd1 vccd1 vccd1 _07222_/A sky130_fd_sc_hd__buf_8
X_09939_ _11665_/Q _09851_/Y _09908_/Y _06969_/X _09938_/Y vssd1 vssd1 vccd1 vccd1
+ _09939_/X sky130_fd_sc_hd__a221o_1
Xfanout863 _05914_/A2 vssd1 vssd1 vccd1 vccd1 _06871_/A2 sky130_fd_sc_hd__buf_6
XFILLER_93_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout874 _10158_/A vssd1 vssd1 vccd1 vccd1 _07939_/A sky130_fd_sc_hd__buf_12
XFILLER_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout885 _06227_/A2 vssd1 vssd1 vccd1 vccd1 _10180_/A sky130_fd_sc_hd__buf_6
XFILLER_19_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout896 _06219_/A2 vssd1 vssd1 vccd1 vccd1 _09359_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_133_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _10021_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11763_ _11763_/CLK _11763_/D vssd1 vssd1 vccd1 vccd1 _11763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10769_/CLK _10714_/D vssd1 vssd1 vccd1 vccd1 _10714_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11765_/CLK _11694_/D vssd1 vssd1 vccd1 vccd1 _11694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10645_ _11270_/CLK _10645_/D vssd1 vssd1 vccd1 vccd1 _10645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10576_ _10769_/CLK _10576_/D vssd1 vssd1 vccd1 vccd1 _10576_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_91_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11644_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _10644_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _11777_/CLK _11128_/D vssd1 vssd1 vccd1 vccd1 _11128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11059_ _11269_/CLK _11059_/D vssd1 vssd1 vccd1 vccd1 _11059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05620_ _05076_/A _11375_/Q _11370_/Q _05620_/B2 _05619_/X vssd1 vssd1 vccd1 vccd1
+ _05621_/B sky130_fd_sc_hd__a221o_4
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05551_ _09552_/A1 _11430_/Q _11424_/Q _11625_/Q vssd1 vssd1 vccd1 vccd1 _05551_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08270_ _10967_/Q _08284_/B vssd1 vssd1 vccd1 vccd1 _08270_/X sky130_fd_sc_hd__or2_1
X_05482_ _10227_/Q input69/X _05508_/S vssd1 vssd1 vccd1 vccd1 _05482_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07221_ _07042_/A _07776_/A2 _07204_/Y _10378_/Q vssd1 vssd1 vccd1 vccd1 _10378_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07152_ _07152_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _09228_/B sky130_fd_sc_hd__nor2_8
X_06103_ _10208_/Q _06351_/A2 _06099_/X _06102_/X vssd1 vssd1 vccd1 vccd1 _06103_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_69_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07083_ _07083_/A _07083_/B vssd1 vssd1 vccd1 vccd1 _07847_/C sky130_fd_sc_hd__nor2_2
XFILLER_106_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06034_ _11562_/Q _09391_/A _06284_/B1 _11552_/Q vssd1 vssd1 vccd1 vccd1 _06034_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07985_ _10817_/Q _07991_/S _07363_/S _07098_/B vssd1 vssd1 vccd1 vccd1 _10817_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09724_ _10350_/Q _09879_/B1 _09882_/B1 _10352_/Q _09723_/X vssd1 vssd1 vccd1 vccd1
+ _09731_/A sky130_fd_sc_hd__a221o_1
XFILLER_80_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06936_ _10213_/Q _06937_/B vssd1 vssd1 vccd1 vccd1 _06938_/B sky130_fd_sc_hd__and2_4
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09655_ _10329_/Q _09570_/A _09566_/D _10335_/Q vssd1 vssd1 vccd1 vccd1 _09655_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06867_ _10250_/Q _06883_/C _06866_/X _06743_/X vssd1 vssd1 vccd1 vccd1 _06868_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08606_ _08793_/A _08606_/B vssd1 vssd1 vccd1 vccd1 _11157_/D sky130_fd_sc_hd__or2_1
X_05818_ _06892_/A _05819_/B vssd1 vssd1 vccd1 vccd1 _05818_/Y sky130_fd_sc_hd__nor2_8
XFILLER_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09586_ _09586_/A _09586_/B _09586_/C _09586_/D vssd1 vssd1 vccd1 vccd1 _09594_/C
+ sky130_fd_sc_hd__nor4_4
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06798_ _11623_/Q _06704_/B _06797_/X vssd1 vssd1 vccd1 vccd1 _10245_/D sky130_fd_sc_hd__a21o_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _08853_/A1 _11118_/Q _08537_/S vssd1 vssd1 vccd1 vccd1 _08538_/B sky130_fd_sc_hd__mux2_1
X_05749_ _05749_/A _05751_/B _05745_/A vssd1 vssd1 vccd1 vccd1 _05749_/X sky130_fd_sc_hd__or3b_4
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08468_ _08749_/A _08468_/B vssd1 vssd1 vccd1 vccd1 _11085_/D sky130_fd_sc_hd__or2_1
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07419_ _10134_/A0 _10486_/Q _07429_/S vssd1 vssd1 vccd1 vccd1 _07420_/B sky130_fd_sc_hd__mux2_1
XFILLER_17_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08399_ _08987_/A1 _08404_/S _08398_/X _08937_/C1 vssd1 vssd1 vccd1 vccd1 _11040_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10430_ _11628_/CLK _10430_/D vssd1 vssd1 vccd1 vccd1 _10430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10361_ _11745_/CLK _10361_/D vssd1 vssd1 vccd1 vccd1 _10361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10292_ _11745_/CLK _10292_/D vssd1 vssd1 vccd1 vccd1 _10292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout660 _11627_/Q vssd1 vssd1 vccd1 vccd1 _05076_/A sky130_fd_sc_hd__buf_12
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout671 _11601_/Q vssd1 vssd1 vccd1 vccd1 _06942_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout682 _05394_/S vssd1 vssd1 vccd1 vccd1 _05432_/S sky130_fd_sc_hd__buf_6
Xfanout693 _05416_/S vssd1 vssd1 vccd1 vccd1 _08956_/B sky130_fd_sc_hd__buf_8
XFILLER_19_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11746_ _11755_/CLK _11746_/D vssd1 vssd1 vccd1 vccd1 _11746_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11677_ _11684_/CLK _11677_/D vssd1 vssd1 vccd1 vccd1 _11677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10628_ _11722_/CLK _10628_/D vssd1 vssd1 vccd1 vccd1 _10628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10559_ _10805_/CLK _10559_/D vssd1 vssd1 vccd1 vccd1 _10559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07770_ _07333_/B _07204_/B _07771_/B1 _10690_/Q _07333_/A vssd1 vssd1 vccd1 vccd1
+ _10690_/D sky130_fd_sc_hd__a221o_1
XFILLER_37_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06721_ _06577_/A _10240_/Q _06855_/B vssd1 vssd1 vccd1 vccd1 _06721_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09440_ _11593_/Q _11652_/Q _09440_/S vssd1 vssd1 vccd1 vccd1 _11593_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06652_ _10387_/Q _07939_/A _08286_/A _10728_/Q vssd1 vssd1 vccd1 vccd1 _06652_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05603_ _05603_/A _05603_/B vssd1 vssd1 vccd1 vccd1 _05603_/Y sky130_fd_sc_hd__nor2_8
XFILLER_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09371_ _11543_/Q _09359_/X _09370_/X vssd1 vssd1 vccd1 vccd1 _11543_/D sky130_fd_sc_hd__a21o_1
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06583_ _10953_/Q _10137_/A _06581_/X _06582_/X vssd1 vssd1 vccd1 vccd1 _06583_/X
+ sky130_fd_sc_hd__o211a_1
X_08322_ _08322_/A _08324_/B vssd1 vssd1 vccd1 vccd1 _08322_/Y sky130_fd_sc_hd__nor2_4
X_05534_ _05630_/A2 _11521_/Q _11518_/Q _05079_/A _05532_/X vssd1 vssd1 vccd1 vccd1
+ _05537_/A sky130_fd_sc_hd__a221o_4
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08253_ _08847_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _10958_/D sky130_fd_sc_hd__or2_1
XFILLER_123_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05465_ _10766_/Q _09879_/A2 _09568_/A _10768_/Q _05460_/X vssd1 vssd1 vccd1 vccd1
+ _05466_/D sky130_fd_sc_hd__a221o_2
X_07204_ _10039_/A _07204_/B vssd1 vssd1 vccd1 vccd1 _07204_/Y sky130_fd_sc_hd__nor2_8
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08184_ _10926_/Q _07052_/A _08197_/S vssd1 vssd1 vccd1 vccd1 _08185_/B sky130_fd_sc_hd__mux2_1
X_05396_ _11210_/Q _11209_/Q _05396_/S vssd1 vssd1 vccd1 vccd1 _05400_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07135_ _10328_/Q _07135_/A2 _07186_/S _07245_/B vssd1 vssd1 vccd1 vccd1 _10328_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07066_ _07211_/A _07074_/S _07065_/X _07141_/B vssd1 vssd1 vccd1 vccd1 _10291_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06017_ _06450_/A _10226_/Q vssd1 vssd1 vccd1 vccd1 _06017_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07968_ _09193_/A _07966_/S _07105_/X vssd1 vssd1 vccd1 vccd1 _07968_/X sky130_fd_sc_hd__a21o_1
XFILLER_87_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06919_ _10153_/A1 _06903_/X _06918_/X _06990_/C1 vssd1 vssd1 vccd1 vccd1 _10200_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09707_ _10407_/Q _09881_/A2 _09876_/B1 _10403_/Q vssd1 vssd1 vccd1 vccd1 _09707_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07899_ _10768_/Q _07901_/B vssd1 vssd1 vccd1 vccd1 _07899_/X sky130_fd_sc_hd__or2_1
XFILLER_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09638_ _11658_/Q _11643_/Q vssd1 vssd1 vccd1 vccd1 _09638_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09569_ _09569_/A _09569_/B _09569_/C _09569_/D vssd1 vssd1 vccd1 vccd1 _09576_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_93_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11600_ _11650_/CLK _11600_/D vssd1 vssd1 vccd1 vccd1 _11600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11531_ _11765_/CLK _11531_/D vssd1 vssd1 vccd1 vccd1 _11531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11462_ _11462_/CLK _11462_/D vssd1 vssd1 vccd1 vccd1 _11462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10413_ _10773_/CLK _10413_/D vssd1 vssd1 vccd1 vccd1 _10413_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11393_ _11393_/CLK _11393_/D vssd1 vssd1 vccd1 vccd1 _11393_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10344_ _10808_/CLK _10344_/D vssd1 vssd1 vccd1 vccd1 _10344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10275_ _11711_/CLK _10275_/D vssd1 vssd1 vccd1 vccd1 _10275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout490 _08843_/C1 vssd1 vssd1 vccd1 vccd1 _07011_/B sky130_fd_sc_hd__buf_6
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11729_ _11762_/CLK _11729_/D vssd1 vssd1 vccd1 vccd1 _11729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05250_ _10982_/Q _10981_/Q _05414_/S vssd1 vssd1 vccd1 vccd1 _05253_/B sky130_fd_sc_hd__mux2_1
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05181_ _10837_/Q _10594_/Q _09538_/A vssd1 vssd1 vccd1 vccd1 _05184_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08940_ input95/X _11329_/Q _08940_/S vssd1 vssd1 vccd1 vccd1 _08941_/B sky130_fd_sc_hd__mux2_1
X_08871_ _08941_/A _08871_/B vssd1 vssd1 vccd1 vccd1 _11292_/D sky130_fd_sc_hd__or2_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07822_ _07048_/A _07839_/A2 _07956_/S _10717_/Q vssd1 vssd1 vccd1 vccd1 _10717_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07753_ _07076_/A _07455_/X _07752_/X _07894_/C1 vssd1 vssd1 vccd1 vccd1 _10677_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06704_ _11618_/Q _06704_/B vssd1 vssd1 vccd1 vccd1 _06704_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07684_ _10640_/Q _07674_/X _07675_/Y _07232_/X vssd1 vssd1 vccd1 vccd1 _10640_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09423_ _11639_/Q _11582_/Q _09704_/B vssd1 vssd1 vccd1 vccd1 _11582_/D sky130_fd_sc_hd__mux2_1
X_06635_ _11134_/Q _06635_/A2 _06635_/B1 _11268_/Q vssd1 vssd1 vccd1 vccd1 _06635_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09354_ _10115_/A0 _11534_/Q _09357_/S vssd1 vssd1 vccd1 vccd1 _11534_/D sky130_fd_sc_hd__mux2_1
X_06566_ _10385_/Q _07939_/A _08286_/A _10726_/Q vssd1 vssd1 vccd1 vccd1 _06566_/X
+ sky130_fd_sc_hd__a22o_1
X_08305_ _10985_/Q _08301_/Y _08304_/Y _08440_/B2 vssd1 vssd1 vccd1 vccd1 _10985_/D
+ sky130_fd_sc_hd__a22o_1
X_05517_ _05626_/A2 _10262_/Q _10257_/Q _05630_/B1 _05516_/X vssd1 vssd1 vccd1 vccd1
+ _05518_/B sky130_fd_sc_hd__a221o_4
X_09285_ _09285_/A1 _09271_/X _09284_/X _09289_/C1 vssd1 vssd1 vccd1 vccd1 _11494_/D
+ sky130_fd_sc_hd__o211a_1
X_06497_ _11148_/Q _07692_/A _06629_/B1 _11099_/Q _07690_/B vssd1 vssd1 vccd1 vccd1
+ _06497_/X sky130_fd_sc_hd__o221a_2
XFILLER_100_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08236_ _10149_/A1 _08325_/B _08235_/X _08753_/C1 vssd1 vssd1 vccd1 vccd1 _10951_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05448_ _10679_/Q _09567_/A _09568_/A _10680_/Q _05435_/X vssd1 vssd1 vccd1 vccd1
+ _05449_/D sky130_fd_sc_hd__a221o_2
XFILLER_14_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08167_ _07048_/A _10909_/Q _08182_/S vssd1 vssd1 vccd1 vccd1 _10909_/D sky130_fd_sc_hd__mux2_1
X_05379_ _05379_/A _05379_/B vssd1 vssd1 vccd1 vccd1 _05379_/Y sky130_fd_sc_hd__nor2_8
XFILLER_118_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07118_ _10315_/Q _07135_/A2 _07186_/S _07052_/X vssd1 vssd1 vccd1 vccd1 _10315_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08098_ _10873_/Q _08902_/B _08362_/B vssd1 vssd1 vccd1 vccd1 _08098_/X sky130_fd_sc_hd__or3_1
XFILLER_109_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07049_ _10280_/Q _07047_/B _07490_/S _07324_/B vssd1 vssd1 vccd1 vccd1 _10280_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_115_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10060_ _11722_/Q _10057_/S _10027_/Y _07040_/B vssd1 vssd1 vccd1 vccd1 _11722_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_102_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10962_ _11575_/CLK _10962_/D vssd1 vssd1 vccd1 vccd1 _10962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10893_ _11601_/CLK _10893_/D vssd1 vssd1 vccd1 vccd1 _10893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11514_ _11763_/CLK _11514_/D vssd1 vssd1 vccd1 vccd1 _11514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ _11473_/CLK _11445_/D vssd1 vssd1 vccd1 vccd1 _11445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11376_ _11495_/CLK _11376_/D vssd1 vssd1 vccd1 vccd1 _11376_/Q sky130_fd_sc_hd__dfxtp_1
X_10327_ _11719_/CLK _10327_/D vssd1 vssd1 vccd1 vccd1 _10327_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _11810_/CLK _10258_/D vssd1 vssd1 vccd1 vccd1 _10258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10189_ _07021_/A _11810_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _11810_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06420_ _07297_/A _06420_/B _06420_/C vssd1 vssd1 vccd1 vccd1 _06420_/X sky130_fd_sc_hd__or3_2
XFILLER_37_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06351_ _10212_/Q _06351_/A2 _06349_/X _06350_/X vssd1 vssd1 vccd1 vccd1 _06351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05302_ _05302_/A _05302_/B vssd1 vssd1 vccd1 vccd1 _05302_/Y sky130_fd_sc_hd__nor2_4
X_09070_ _09141_/A1 _09060_/X _09069_/X _09168_/C1 vssd1 vssd1 vccd1 vccd1 _11383_/D
+ sky130_fd_sc_hd__o211a_1
X_06282_ _11516_/Q _09314_/A _06278_/X _06281_/X vssd1 vssd1 vccd1 vccd1 _06282_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ _10835_/Q _08037_/B vssd1 vssd1 vccd1 vccd1 _08021_/X sky130_fd_sc_hd__or2_1
X_05233_ _09539_/A _10950_/Q _05225_/X _05228_/X _05229_/X vssd1 vssd1 vccd1 vccd1
+ _05233_/X sky130_fd_sc_hd__a2111o_1
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05164_ _10597_/Q _11077_/Q _05394_/S vssd1 vssd1 vccd1 vccd1 _05167_/B sky130_fd_sc_hd__mux2_1
XFILLER_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09972_ _08092_/A _11672_/Q _09975_/S vssd1 vssd1 vccd1 vccd1 _11672_/D sky130_fd_sc_hd__mux2_1
X_05095_ _11871_/A vssd1 vssd1 vccd1 vccd1 _05095_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08923_ _08987_/A1 _08940_/S _08922_/X _08943_/C1 vssd1 vssd1 vccd1 vccd1 _11320_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08854_ _08855_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08894_/B sky130_fd_sc_hd__nor2_4
XFILLER_44_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07805_ _07028_/A _10710_/Q _09193_/B vssd1 vssd1 vccd1 vccd1 _07806_/B sky130_fd_sc_hd__mux2_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08785_ _08875_/A _08785_/B vssd1 vssd1 vccd1 vccd1 _11248_/D sky130_fd_sc_hd__or2_1
X_05997_ _10912_/Q _06591_/A2 _05865_/B _11769_/Q vssd1 vssd1 vccd1 vccd1 _05997_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_73_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ _10669_/Q _07750_/B vssd1 vssd1 vccd1 vccd1 _07736_/X sky130_fd_sc_hd__or2_1
XFILLER_38_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07667_ _10628_/Q _07665_/S _07249_/S _07141_/X vssd1 vssd1 vccd1 vccd1 _10628_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06618_ _11871_/A _06612_/X _06617_/X _06576_/A vssd1 vssd1 vccd1 vccd1 _06618_/X
+ sky130_fd_sc_hd__a31o_1
X_09406_ _09681_/B _09406_/B vssd1 vssd1 vccd1 vccd1 _09407_/B sky130_fd_sc_hd__nor2_8
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07598_ _09206_/A _08850_/S vssd1 vssd1 vccd1 vccd1 _07598_/Y sky130_fd_sc_hd__nand2_2
XFILLER_41_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09337_ _10171_/A1 _09343_/B _08851_/A vssd1 vssd1 vccd1 vccd1 _09337_/X sky130_fd_sc_hd__a21o_1
X_06549_ _10922_/Q _06591_/A2 _06126_/B _11218_/Q vssd1 vssd1 vccd1 vccd1 _06552_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09268_ _10106_/A1 _09266_/B _08761_/A vssd1 vssd1 vccd1 vccd1 _09268_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08219_ _08970_/A1 _10944_/Q _08219_/S vssd1 vssd1 vccd1 vccd1 _08220_/B sky130_fd_sc_hd__mux2_1
XFILLER_153_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09199_ _07143_/X _09192_/B _09190_/Y _11446_/Q _09192_/A vssd1 vssd1 vccd1 vccd1
+ _11446_/D sky130_fd_sc_hd__a221o_1
XFILLER_101_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _11629_/CLK _11230_/D vssd1 vssd1 vccd1 vccd1 _11230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _11332_/CLK _11161_/D vssd1 vssd1 vccd1 vccd1 _11161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10112_ _10112_/A0 _11759_/Q _10118_/S vssd1 vssd1 vccd1 vccd1 _11759_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11092_ _11312_/CLK _11092_/D vssd1 vssd1 vccd1 vccd1 _11092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10043_ _10043_/A _10043_/B vssd1 vssd1 vccd1 vccd1 _11712_/D sky130_fd_sc_hd__or2_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10945_ _11023_/CLK _10945_/D vssd1 vssd1 vccd1 vccd1 _10945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_45_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _11755_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10876_ _10932_/CLK _10876_/D vssd1 vssd1 vccd1 vccd1 _10876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_4 _05313_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11428_ _11428_/CLK _11428_/D vssd1 vssd1 vccd1 vccd1 _11428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ _11809_/CLK _11359_/D vssd1 vssd1 vccd1 vccd1 _11359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05920_ _11035_/Q _08383_/A _08245_/A _10957_/Q vssd1 vssd1 vccd1 vccd1 _05922_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1060 _10166_/A1 vssd1 vssd1 vccd1 vccd1 _09090_/A1 sky130_fd_sc_hd__buf_6
Xfanout1071 input110/X vssd1 vssd1 vccd1 vccd1 _10142_/A1 sky130_fd_sc_hd__buf_12
XFILLER_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05851_ _11452_/Q _06799_/A2 _06999_/A _10339_/Q _06651_/C1 vssd1 vssd1 vccd1 vccd1
+ _05851_/X sky130_fd_sc_hd__o221a_1
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08570_ _08749_/A _08570_/B vssd1 vssd1 vccd1 vccd1 _11139_/D sky130_fd_sc_hd__or2_1
X_05782_ _10746_/Q _07853_/A _07152_/A _10338_/Q _05781_/X vssd1 vssd1 vccd1 vccd1
+ _05782_/X sky130_fd_sc_hd__o221a_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07521_ _07025_/A _10545_/Q _07533_/S vssd1 vssd1 vccd1 vccd1 _07522_/B sky130_fd_sc_hd__mux2_1
XFILLER_78_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07452_ _10503_/Q _07441_/Y _07443_/Y _07451_/X vssd1 vssd1 vccd1 vccd1 _10503_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06403_ _06397_/X _06402_/X _11870_/A vssd1 vssd1 vccd1 vccd1 _06403_/X sky130_fd_sc_hd__o21a_1
X_07383_ _08733_/A _07383_/B vssd1 vssd1 vccd1 vccd1 _10466_/D sky130_fd_sc_hd__or2_1
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09122_ _09283_/A1 _09110_/X _09121_/X _09122_/C1 vssd1 vssd1 vccd1 vccd1 _11407_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06334_ _10447_/Q _07222_/A _07819_/A _10304_/Q vssd1 vssd1 vccd1 vccd1 _06334_/X
+ sky130_fd_sc_hd__o22a_1
X_09053_ _10023_/A0 _09055_/B _09129_/B1 vssd1 vssd1 vccd1 vccd1 _09053_/X sky130_fd_sc_hd__a21o_1
XFILLER_135_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06265_ _10640_/Q _06538_/B1 _06264_/X _06265_/C1 vssd1 vssd1 vccd1 vccd1 _06265_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08004_ _08839_/A _08004_/B vssd1 vssd1 vccd1 vccd1 _10826_/D sky130_fd_sc_hd__or2_1
X_05216_ _05426_/S _11059_/Q _10854_/Q _09681_/A _05215_/X vssd1 vssd1 vccd1 vccd1
+ _05224_/A sky130_fd_sc_hd__a221o_2
XFILLER_135_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06196_ _10480_/Q _06803_/A2 _06685_/B _11701_/Q vssd1 vssd1 vccd1 vccd1 _06196_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_102_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05147_ _10944_/Q _10943_/Q _05430_/S vssd1 vssd1 vccd1 vccd1 _05151_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05078_ _05078_/A vssd1 vssd1 vccd1 vccd1 _05078_/Y sky130_fd_sc_hd__clkinv_2
X_09955_ _09955_/A _09955_/B _09955_/C _09955_/D vssd1 vssd1 vccd1 vccd1 _09958_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08906_ _08907_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08906_/Y sky130_fd_sc_hd__nor2_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _10557_/Q _09886_/A2 _09886_/B1 _10579_/Q _09871_/X vssd1 vssd1 vccd1 vccd1
+ _09887_/D sky130_fd_sc_hd__a221o_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _07107_/A _08838_/S _08836_/X _08841_/C1 vssd1 vssd1 vccd1 vccd1 _11276_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapped_tms1x00_1103 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1103/HI io_oeb[33] sky130_fd_sc_hd__conb_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1114 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_1114/HI io_out[6] sky130_fd_sc_hd__conb_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_tms1x00_1125 vssd1 vssd1 vccd1 vccd1 io_oeb[2] wrapped_tms1x00_1125/LO sky130_fd_sc_hd__conb_1
X_08768_ _09275_/A1 _11240_/Q _08802_/S vssd1 vssd1 vccd1 vccd1 _08769_/B sky130_fd_sc_hd__mux2_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07719_ _10023_/A0 _07755_/A2 _07718_/X _07868_/C1 vssd1 vssd1 vccd1 vccd1 _10660_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _11204_/Q _08705_/B vssd1 vssd1 vccd1 vccd1 _08699_/X sky130_fd_sc_hd__or2_1
XFILLER_92_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10730_ _11711_/CLK _10730_/D vssd1 vssd1 vccd1 vccd1 _10730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10661_ _11465_/CLK _10661_/D vssd1 vssd1 vccd1 vccd1 _10661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10592_ _11657_/CLK _10592_/D vssd1 vssd1 vccd1 vccd1 _10592_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11213_ _11220_/CLK _11213_/D vssd1 vssd1 vccd1 vccd1 _11213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11144_ _11652_/CLK _11144_/D vssd1 vssd1 vccd1 vccd1 _11144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11075_ _11177_/CLK _11075_/D vssd1 vssd1 vccd1 vccd1 _11075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10026_ _10026_/A _10026_/B vssd1 vssd1 vccd1 vccd1 _11703_/D sky130_fd_sc_hd__or2_1
XFILLER_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10928_ _10932_/CLK _10928_/D vssd1 vssd1 vccd1 vccd1 _10928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ _10939_/CLK _10859_/D vssd1 vssd1 vccd1 vccd1 _10859_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06050_ _11317_/Q _06413_/A2 _06455_/B1 _11243_/Q vssd1 vssd1 vccd1 vccd1 _06050_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout308 _07455_/X vssd1 vssd1 vccd1 vccd1 _07755_/A2 sky130_fd_sc_hd__buf_6
Xfanout319 _07337_/X vssd1 vssd1 vccd1 vccd1 _07350_/S sky130_fd_sc_hd__buf_6
XFILLER_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09740_ _09908_/A _09740_/B vssd1 vssd1 vccd1 vccd1 _09740_/Y sky130_fd_sc_hd__nor2_2
X_06952_ _10218_/Q _06951_/X _09416_/A vssd1 vssd1 vccd1 vccd1 _10218_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
.ends

