// This is the unpowered netlist.
module wrapped_tms1x00 (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out,
    oram_addr,
    oram_value);
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [8:0] oram_addr;
 input [31:0] oram_value;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire net93;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net94;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net95;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire clknet_0_wb_clk_i;
 wire net96;
 wire net97;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net59;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net60;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net61;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net92;
 wire \tms1x00.CL ;
 wire \tms1x00.PA[0] ;
 wire \tms1x00.PA[1] ;
 wire \tms1x00.PA[2] ;
 wire \tms1x00.PA[3] ;
 wire \tms1x00.PB[0] ;
 wire \tms1x00.PB[1] ;
 wire \tms1x00.PB[2] ;
 wire \tms1x00.PB[3] ;
 wire \tms1x00.PC[0] ;
 wire \tms1x00.PC[1] ;
 wire \tms1x00.PC[2] ;
 wire \tms1x00.PC[3] ;
 wire \tms1x00.PC[4] ;
 wire \tms1x00.PC[5] ;
 wire \tms1x00.SR[0] ;
 wire \tms1x00.SR[1] ;
 wire \tms1x00.SR[2] ;
 wire \tms1x00.SR[3] ;
 wire \tms1x00.SR[4] ;
 wire \tms1x00.SR[5] ;
 wire \tms1x00.ins_in[0] ;
 wire \tms1x00.ins_in[1] ;
 wire \tms1x00.ins_in[2] ;
 wire \tms1x00.ins_in[3] ;
 wire \tms1x00.ins_in[4] ;
 wire \tms1x00.ins_in[5] ;
 wire \tms1x00.ins_in[6] ;
 wire \tms1x00.ins_in[7] ;
 wire \tms1x00.rom_addr[0] ;
 wire \tms1x00.rom_addr[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;

 sky130_fd_sc_hd__buf_2 _156_ (.A(net12),
    .X(_044_));
 sky130_fd_sc_hd__buf_2 _157_ (.A(_044_),
    .X(_045_));
 sky130_fd_sc_hd__nor2_1 _158_ (.A(_045_),
    .B(net14),
    .Y(_000_));
 sky130_fd_sc_hd__nor2_1 _159_ (.A(net15),
    .B(net14),
    .Y(_046_));
 sky130_fd_sc_hd__and3b_1 _160_ (.A_N(net15),
    .B(net14),
    .C(net16),
    .X(_047_));
 sky130_fd_sc_hd__or3_1 _161_ (.A(net12),
    .B(_046_),
    .C(_047_),
    .X(_048_));
 sky130_fd_sc_hd__nand2_1 _162_ (.A(net15),
    .B(net14),
    .Y(_049_));
 sky130_fd_sc_hd__and2b_1 _163_ (.A_N(_048_),
    .B(_049_),
    .X(_050_));
 sky130_fd_sc_hd__clkbuf_1 _164_ (.A(_050_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _165_ (.A0(_049_),
    .A1(net14),
    .S(net16),
    .X(_051_));
 sky130_fd_sc_hd__nor2_1 _166_ (.A(_045_),
    .B(_051_),
    .Y(_002_));
 sky130_fd_sc_hd__and2_2 _167_ (.A(net16),
    .B(_046_),
    .X(_052_));
 sky130_fd_sc_hd__or2_1 _168_ (.A(net12),
    .B(_052_),
    .X(_053_));
 sky130_fd_sc_hd__buf_2 _169_ (.A(_053_),
    .X(_054_));
 sky130_fd_sc_hd__nand2_1 _170_ (.A(net16),
    .B(_046_),
    .Y(_055_));
 sky130_fd_sc_hd__or2_1 _171_ (.A(_044_),
    .B(_055_),
    .X(_056_));
 sky130_fd_sc_hd__clkbuf_4 _172_ (.A(\tms1x00.rom_addr[1] ),
    .X(_057_));
 sky130_fd_sc_hd__mux4_2 _173_ (.A0(net1),
    .A1(net3),
    .A2(net4),
    .A3(net5),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_057_),
    .X(_058_));
 sky130_fd_sc_hd__o22a_1 _174_ (.A1(\tms1x00.ins_in[0] ),
    .A2(_054_),
    .B1(_056_),
    .B2(_058_),
    .X(_003_));
 sky130_fd_sc_hd__mux4_2 _175_ (.A0(net3),
    .A1(net4),
    .A2(net5),
    .A3(net6),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_057_),
    .X(_059_));
 sky130_fd_sc_hd__o22a_1 _176_ (.A1(\tms1x00.ins_in[1] ),
    .A2(_054_),
    .B1(_056_),
    .B2(_059_),
    .X(_004_));
 sky130_fd_sc_hd__nor2_1 _177_ (.A(_044_),
    .B(_055_),
    .Y(_060_));
 sky130_fd_sc_hd__mux2_1 _178_ (.A0(net4),
    .A1(net5),
    .S(\tms1x00.rom_addr[0] ),
    .X(_061_));
 sky130_fd_sc_hd__or2_1 _179_ (.A(_057_),
    .B(_061_),
    .X(_062_));
 sky130_fd_sc_hd__mux2_1 _180_ (.A0(net6),
    .A1(net7),
    .S(\tms1x00.rom_addr[0] ),
    .X(_063_));
 sky130_fd_sc_hd__or2b_1 _181_ (.A(_063_),
    .B_N(_057_),
    .X(_064_));
 sky130_fd_sc_hd__nor2_1 _182_ (.A(_044_),
    .B(_052_),
    .Y(_065_));
 sky130_fd_sc_hd__a32o_1 _183_ (.A1(_060_),
    .A2(_062_),
    .A3(_064_),
    .B1(_065_),
    .B2(\tms1x00.ins_in[2] ),
    .X(_005_));
 sky130_fd_sc_hd__mux4_2 _184_ (.A0(net5),
    .A1(net6),
    .A2(net7),
    .A3(net8),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_057_),
    .X(_066_));
 sky130_fd_sc_hd__o21ba_1 _185_ (.A1(\tms1x00.ins_in[3] ),
    .A2(_052_),
    .B1_N(_044_),
    .X(_067_));
 sky130_fd_sc_hd__o21a_1 _186_ (.A1(_055_),
    .A2(_066_),
    .B1(_067_),
    .X(_006_));
 sky130_fd_sc_hd__or2_1 _187_ (.A(_057_),
    .B(_063_),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _188_ (.A0(net8),
    .A1(net9),
    .S(\tms1x00.rom_addr[0] ),
    .X(_069_));
 sky130_fd_sc_hd__or2b_1 _189_ (.A(_069_),
    .B_N(_057_),
    .X(_070_));
 sky130_fd_sc_hd__a32o_1 _190_ (.A1(_060_),
    .A2(_068_),
    .A3(_070_),
    .B1(_065_),
    .B2(\tms1x00.ins_in[4] ),
    .X(_007_));
 sky130_fd_sc_hd__mux4_2 _191_ (.A0(net7),
    .A1(net8),
    .A2(net9),
    .A3(net10),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_071_));
 sky130_fd_sc_hd__mux2_1 _192_ (.A0(\tms1x00.ins_in[5] ),
    .A1(_071_),
    .S(_052_),
    .X(_072_));
 sky130_fd_sc_hd__or2_1 _193_ (.A(_045_),
    .B(_072_),
    .X(_073_));
 sky130_fd_sc_hd__clkbuf_1 _194_ (.A(_073_),
    .X(_008_));
 sky130_fd_sc_hd__mux4_2 _195_ (.A0(net8),
    .A1(net9),
    .A2(net10),
    .A3(net11),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_057_),
    .X(_074_));
 sky130_fd_sc_hd__a22o_1 _196_ (.A1(\tms1x00.ins_in[6] ),
    .A2(_065_),
    .B1(_060_),
    .B2(_074_),
    .X(_009_));
 sky130_fd_sc_hd__mux4_2 _197_ (.A0(net9),
    .A1(net10),
    .A2(net11),
    .A3(net2),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_057_),
    .X(_075_));
 sky130_fd_sc_hd__a22o_1 _198_ (.A1(\tms1x00.ins_in[7] ),
    .A2(_065_),
    .B1(_060_),
    .B2(_075_),
    .X(_010_));
 sky130_fd_sc_hd__clkinv_2 _199_ (.A(net13),
    .Y(_076_));
 sky130_fd_sc_hd__or2_1 _200_ (.A(net16),
    .B(_049_),
    .X(_077_));
 sky130_fd_sc_hd__or4_1 _201_ (.A(\tms1x00.ins_in[3] ),
    .B(\tms1x00.ins_in[2] ),
    .C(\tms1x00.ins_in[1] ),
    .D(\tms1x00.ins_in[0] ),
    .X(_078_));
 sky130_fd_sc_hd__nand2_1 _202_ (.A(\tms1x00.ins_in[6] ),
    .B(\tms1x00.ins_in[4] ),
    .Y(_079_));
 sky130_fd_sc_hd__or4_1 _203_ (.A(\tms1x00.ins_in[5] ),
    .B(_077_),
    .C(_078_),
    .D(_079_),
    .X(_080_));
 sky130_fd_sc_hd__mux2_1 _204_ (.A0(\tms1x00.ins_in[7] ),
    .A1(_076_),
    .S(_080_),
    .X(_081_));
 sky130_fd_sc_hd__nor2_1 _205_ (.A(_045_),
    .B(_081_),
    .Y(_011_));
 sky130_fd_sc_hd__and4b_1 _206_ (.A_N(net15),
    .B(net14),
    .C(\tms1x00.ins_in[0] ),
    .D(net16),
    .X(_082_));
 sky130_fd_sc_hd__buf_2 _207_ (.A(_082_),
    .X(_083_));
 sky130_fd_sc_hd__and2_2 _208_ (.A(\tms1x00.ins_in[1] ),
    .B(_083_),
    .X(_084_));
 sky130_fd_sc_hd__nor4_1 _209_ (.A(\tms1x00.ins_in[3] ),
    .B(\tms1x00.ins_in[2] ),
    .C(\tms1x00.ins_in[1] ),
    .D(\tms1x00.ins_in[0] ),
    .Y(_085_));
 sky130_fd_sc_hd__and4_1 _210_ (.A(\tms1x00.ins_in[7] ),
    .B(\tms1x00.ins_in[6] ),
    .C(\tms1x00.ins_in[5] ),
    .D(\tms1x00.ins_in[4] ),
    .X(_086_));
 sky130_fd_sc_hd__and4_1 _211_ (.A(\tms1x00.CL ),
    .B(_047_),
    .C(_085_),
    .D(_086_),
    .X(_087_));
 sky130_fd_sc_hd__buf_2 _212_ (.A(_087_),
    .X(_088_));
 sky130_fd_sc_hd__nor2_1 _213_ (.A(_045_),
    .B(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__o21a_1 _214_ (.A1(\tms1x00.CL ),
    .A2(_084_),
    .B1(_089_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _215_ (.A0(\tms1x00.PB[0] ),
    .A1(\tms1x00.PA[0] ),
    .S(_084_),
    .X(_090_));
 sky130_fd_sc_hd__or4b_1 _216_ (.A(\tms1x00.ins_in[2] ),
    .B(\tms1x00.ins_in[1] ),
    .C(\tms1x00.ins_in[0] ),
    .D_N(\tms1x00.ins_in[3] ),
    .X(_091_));
 sky130_fd_sc_hd__or2_2 _217_ (.A(_077_),
    .B(_091_),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _218_ (.A0(\tms1x00.ins_in[4] ),
    .A1(_090_),
    .S(_092_),
    .X(_093_));
 sky130_fd_sc_hd__or2_1 _219_ (.A(_045_),
    .B(_093_),
    .X(_094_));
 sky130_fd_sc_hd__clkbuf_1 _220_ (.A(_094_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _221_ (.A0(\tms1x00.PB[1] ),
    .A1(\tms1x00.PA[1] ),
    .S(_084_),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _222_ (.A0(\tms1x00.ins_in[5] ),
    .A1(_095_),
    .S(_092_),
    .X(_096_));
 sky130_fd_sc_hd__or2_1 _223_ (.A(_045_),
    .B(_096_),
    .X(_097_));
 sky130_fd_sc_hd__clkbuf_1 _224_ (.A(_097_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _225_ (.A0(\tms1x00.PB[2] ),
    .A1(\tms1x00.PA[2] ),
    .S(_084_),
    .X(_098_));
 sky130_fd_sc_hd__mux2_1 _226_ (.A0(\tms1x00.ins_in[6] ),
    .A1(_098_),
    .S(_092_),
    .X(_099_));
 sky130_fd_sc_hd__or2_1 _227_ (.A(_045_),
    .B(_099_),
    .X(_100_));
 sky130_fd_sc_hd__clkbuf_1 _228_ (.A(_100_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _229_ (.A0(\tms1x00.PB[3] ),
    .A1(\tms1x00.PA[3] ),
    .S(_084_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _230_ (.A0(\tms1x00.ins_in[7] ),
    .A1(_101_),
    .S(_092_),
    .X(_102_));
 sky130_fd_sc_hd__or2_1 _231_ (.A(_044_),
    .B(_102_),
    .X(_103_));
 sky130_fd_sc_hd__clkbuf_1 _232_ (.A(_103_),
    .X(_016_));
 sky130_fd_sc_hd__inv_2 _233_ (.A(\tms1x00.ins_in[1] ),
    .Y(_104_));
 sky130_fd_sc_hd__or2b_1 _234_ (.A(\tms1x00.CL ),
    .B_N(\tms1x00.ins_in[0] ),
    .X(_105_));
 sky130_fd_sc_hd__or4b_4 _235_ (.A(_104_),
    .B(_105_),
    .C(net12),
    .D_N(_047_),
    .X(_106_));
 sky130_fd_sc_hd__mux2_1 _236_ (.A0(\tms1x00.PC[0] ),
    .A1(\tms1x00.SR[0] ),
    .S(_106_),
    .X(_107_));
 sky130_fd_sc_hd__clkbuf_1 _237_ (.A(_107_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _238_ (.A0(\tms1x00.PC[1] ),
    .A1(\tms1x00.SR[1] ),
    .S(_106_),
    .X(_108_));
 sky130_fd_sc_hd__clkbuf_1 _239_ (.A(_108_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _240_ (.A0(\tms1x00.PC[2] ),
    .A1(\tms1x00.SR[2] ),
    .S(_106_),
    .X(_109_));
 sky130_fd_sc_hd__clkbuf_1 _241_ (.A(_109_),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _242_ (.A0(\tms1x00.PC[3] ),
    .A1(\tms1x00.SR[3] ),
    .S(_106_),
    .X(_110_));
 sky130_fd_sc_hd__clkbuf_1 _243_ (.A(_110_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _244_ (.A0(\tms1x00.PC[4] ),
    .A1(\tms1x00.SR[4] ),
    .S(_106_),
    .X(_111_));
 sky130_fd_sc_hd__clkbuf_1 _245_ (.A(_111_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _246_ (.A0(\tms1x00.PC[5] ),
    .A1(\tms1x00.SR[5] ),
    .S(_106_),
    .X(_112_));
 sky130_fd_sc_hd__clkbuf_1 _247_ (.A(_112_),
    .X(_022_));
 sky130_fd_sc_hd__or3_1 _248_ (.A(\tms1x00.PC[0] ),
    .B(_083_),
    .C(_088_),
    .X(_113_));
 sky130_fd_sc_hd__and2b_1 _249_ (.A_N(\tms1x00.ins_in[2] ),
    .B(_083_),
    .X(_114_));
 sky130_fd_sc_hd__and3_1 _250_ (.A(\tms1x00.CL ),
    .B(_085_),
    .C(_086_),
    .X(_115_));
 sky130_fd_sc_hd__a2bb2o_1 _251_ (.A1_N(_088_),
    .A2_N(_114_),
    .B1(\tms1x00.SR[0] ),
    .B2(_115_),
    .X(_116_));
 sky130_fd_sc_hd__and3_1 _252_ (.A(_052_),
    .B(_113_),
    .C(_116_),
    .X(_117_));
 sky130_fd_sc_hd__a21oi_1 _253_ (.A1(_113_),
    .A2(_116_),
    .B1(_052_),
    .Y(_118_));
 sky130_fd_sc_hd__nor3_1 _254_ (.A(_045_),
    .B(_117_),
    .C(_118_),
    .Y(_023_));
 sky130_fd_sc_hd__nor2_2 _255_ (.A(_083_),
    .B(_088_),
    .Y(_119_));
 sky130_fd_sc_hd__a22o_1 _256_ (.A1(\tms1x00.ins_in[3] ),
    .A2(_083_),
    .B1(_088_),
    .B2(\tms1x00.SR[1] ),
    .X(_120_));
 sky130_fd_sc_hd__a21oi_1 _257_ (.A1(\tms1x00.PC[1] ),
    .A2(_119_),
    .B1(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__nor2_1 _258_ (.A(_054_),
    .B(_121_),
    .Y(_024_));
 sky130_fd_sc_hd__a22o_1 _259_ (.A1(\tms1x00.ins_in[4] ),
    .A2(_083_),
    .B1(_088_),
    .B2(\tms1x00.SR[2] ),
    .X(_122_));
 sky130_fd_sc_hd__a21oi_1 _260_ (.A1(\tms1x00.PC[2] ),
    .A2(_119_),
    .B1(_122_),
    .Y(_123_));
 sky130_fd_sc_hd__nor2_1 _261_ (.A(_054_),
    .B(_123_),
    .Y(_025_));
 sky130_fd_sc_hd__a22o_1 _262_ (.A1(\tms1x00.ins_in[5] ),
    .A2(_083_),
    .B1(_088_),
    .B2(\tms1x00.SR[3] ),
    .X(_124_));
 sky130_fd_sc_hd__a21oi_1 _263_ (.A1(\tms1x00.PC[3] ),
    .A2(_119_),
    .B1(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__nor2_1 _264_ (.A(_054_),
    .B(_125_),
    .Y(_026_));
 sky130_fd_sc_hd__a22o_1 _265_ (.A1(\tms1x00.ins_in[6] ),
    .A2(_083_),
    .B1(_088_),
    .B2(\tms1x00.SR[4] ),
    .X(_126_));
 sky130_fd_sc_hd__a21oi_1 _266_ (.A1(\tms1x00.PC[4] ),
    .A2(_119_),
    .B1(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__nor2_1 _267_ (.A(_054_),
    .B(_127_),
    .Y(_027_));
 sky130_fd_sc_hd__a22o_1 _268_ (.A1(\tms1x00.ins_in[7] ),
    .A2(_083_),
    .B1(_088_),
    .B2(\tms1x00.SR[5] ),
    .X(_128_));
 sky130_fd_sc_hd__a21oi_1 _269_ (.A1(\tms1x00.PC[5] ),
    .A2(_119_),
    .B1(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__nor2_1 _270_ (.A(_054_),
    .B(_129_),
    .Y(_028_));
 sky130_fd_sc_hd__or3_1 _271_ (.A(net12),
    .B(net16),
    .C(net15),
    .X(_130_));
 sky130_fd_sc_hd__clkbuf_4 _272_ (.A(_130_),
    .X(_131_));
 sky130_fd_sc_hd__mux2_1 _273_ (.A0(\tms1x00.PC[0] ),
    .A1(\tms1x00.rom_addr[0] ),
    .S(_131_),
    .X(_132_));
 sky130_fd_sc_hd__clkbuf_1 _274_ (.A(_132_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _275_ (.A0(\tms1x00.PC[1] ),
    .A1(_057_),
    .S(_131_),
    .X(_133_));
 sky130_fd_sc_hd__clkbuf_1 _276_ (.A(_133_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _277_ (.A0(\tms1x00.PC[2] ),
    .A1(net18),
    .S(_131_),
    .X(_134_));
 sky130_fd_sc_hd__clkbuf_1 _278_ (.A(_134_),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _279_ (.A0(\tms1x00.PC[3] ),
    .A1(net19),
    .S(_131_),
    .X(_135_));
 sky130_fd_sc_hd__clkbuf_1 _280_ (.A(_135_),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _281_ (.A0(\tms1x00.PC[4] ),
    .A1(net20),
    .S(_131_),
    .X(_136_));
 sky130_fd_sc_hd__clkbuf_1 _282_ (.A(_136_),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _283_ (.A0(\tms1x00.PC[5] ),
    .A1(net21),
    .S(_131_),
    .X(_137_));
 sky130_fd_sc_hd__clkbuf_1 _284_ (.A(_137_),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _285_ (.A0(\tms1x00.PA[0] ),
    .A1(net22),
    .S(_131_),
    .X(_138_));
 sky130_fd_sc_hd__clkbuf_1 _286_ (.A(_138_),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _287_ (.A0(\tms1x00.PA[1] ),
    .A1(net23),
    .S(_131_),
    .X(_139_));
 sky130_fd_sc_hd__clkbuf_1 _288_ (.A(_139_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _289_ (.A0(\tms1x00.PA[2] ),
    .A1(net24),
    .S(_131_),
    .X(_140_));
 sky130_fd_sc_hd__clkbuf_1 _290_ (.A(_140_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _291_ (.A0(\tms1x00.PA[3] ),
    .A1(net25),
    .S(_131_),
    .X(_141_));
 sky130_fd_sc_hd__clkbuf_1 _292_ (.A(_141_),
    .X(_038_));
 sky130_fd_sc_hd__nand2_1 _293_ (.A(\tms1x00.ins_in[5] ),
    .B(\tms1x00.ins_in[4] ),
    .Y(_142_));
 sky130_fd_sc_hd__or4_1 _294_ (.A(\tms1x00.ins_in[6] ),
    .B(_077_),
    .C(_078_),
    .D(_142_),
    .X(_143_));
 sky130_fd_sc_hd__mux2_1 _295_ (.A0(\tms1x00.ins_in[7] ),
    .A1(net17),
    .S(_143_),
    .X(_144_));
 sky130_fd_sc_hd__and2b_1 _296_ (.A_N(_045_),
    .B(_144_),
    .X(_145_));
 sky130_fd_sc_hd__clkbuf_1 _297_ (.A(_145_),
    .X(_039_));
 sky130_fd_sc_hd__nand2_1 _298_ (.A(_085_),
    .B(_086_),
    .Y(_146_));
 sky130_fd_sc_hd__a21boi_4 _299_ (.A1(_146_),
    .A2(_105_),
    .B1_N(_047_),
    .Y(_147_));
 sky130_fd_sc_hd__mux2_1 _300_ (.A0(\tms1x00.PA[3] ),
    .A1(\tms1x00.PB[3] ),
    .S(_147_),
    .X(_148_));
 sky130_fd_sc_hd__or2_1 _301_ (.A(_044_),
    .B(_148_),
    .X(_149_));
 sky130_fd_sc_hd__clkbuf_1 _302_ (.A(_149_),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _303_ (.A0(\tms1x00.PA[2] ),
    .A1(\tms1x00.PB[2] ),
    .S(_147_),
    .X(_150_));
 sky130_fd_sc_hd__or2_1 _304_ (.A(_044_),
    .B(_150_),
    .X(_151_));
 sky130_fd_sc_hd__clkbuf_1 _305_ (.A(_151_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _306_ (.A0(\tms1x00.PA[1] ),
    .A1(\tms1x00.PB[1] ),
    .S(_147_),
    .X(_152_));
 sky130_fd_sc_hd__or2_1 _307_ (.A(_044_),
    .B(_152_),
    .X(_153_));
 sky130_fd_sc_hd__clkbuf_1 _308_ (.A(_153_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _309_ (.A0(\tms1x00.PA[0] ),
    .A1(\tms1x00.PB[0] ),
    .S(_147_),
    .X(_154_));
 sky130_fd_sc_hd__or2_1 _310_ (.A(_044_),
    .B(_154_),
    .X(_155_));
 sky130_fd_sc_hd__clkbuf_1 _311_ (.A(_155_),
    .X(_043_));
 sky130_fd_sc_hd__dfxtp_4 _312_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_000_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_4 _313_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_001_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_4 _314_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_002_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _315_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_003_),
    .Q(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__dfxtp_2 _316_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_004_),
    .Q(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _317_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_005_),
    .Q(\tms1x00.ins_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _318_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_006_),
    .Q(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__dfxtp_2 _319_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_007_),
    .Q(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _320_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_008_),
    .Q(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__dfxtp_2 _321_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_009_),
    .Q(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__dfxtp_2 _322_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_010_),
    .Q(\tms1x00.ins_in[7] ));
 sky130_fd_sc_hd__dfxtp_4 _323_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_011_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _324_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_012_),
    .Q(\tms1x00.CL ));
 sky130_fd_sc_hd__dfxtp_1 _325_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_013_),
    .Q(\tms1x00.PB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _326_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_014_),
    .Q(\tms1x00.PB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _327_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_015_),
    .Q(\tms1x00.PB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _328_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_016_),
    .Q(\tms1x00.PB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _329_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_017_),
    .Q(\tms1x00.SR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _330_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_018_),
    .Q(\tms1x00.SR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _331_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_019_),
    .Q(\tms1x00.SR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _332_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_020_),
    .Q(\tms1x00.SR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _333_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_021_),
    .Q(\tms1x00.SR[4] ));
 sky130_fd_sc_hd__dfxtp_1 _334_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_022_),
    .Q(\tms1x00.SR[5] ));
 sky130_fd_sc_hd__dfxtp_1 _335_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_023_),
    .Q(\tms1x00.PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _336_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_024_),
    .Q(\tms1x00.PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _337_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_025_),
    .Q(\tms1x00.PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _338_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_026_),
    .Q(\tms1x00.PC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _339_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_027_),
    .Q(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _340_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_028_),
    .Q(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__dfxtp_4 _341_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_029_),
    .Q(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _342_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_030_),
    .Q(\tms1x00.rom_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _343_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_031_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _344_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_032_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _345_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_033_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _346_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_034_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_2 _347_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_035_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_2 _348_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_036_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_2 _349_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_037_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_2 _350_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_038_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_4 _351_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_039_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _352_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_040_),
    .Q(\tms1x00.PA[3] ));
 sky130_fd_sc_hd__dfxtp_1 _353_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_041_),
    .Q(\tms1x00.PA[2] ));
 sky130_fd_sc_hd__dfxtp_1 _354_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_042_),
    .Q(\tms1x00.PA[1] ));
 sky130_fd_sc_hd__dfxtp_1 _355_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_043_),
    .Q(\tms1x00.PA[0] ));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_93 (.HI(net93));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_94 (.HI(net94));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_95 (.HI(net95));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_96 (.HI(net96));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_97 (.HI(net97));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_92 (.HI(net92));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(oram_value[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(oram_value[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(oram_value[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(oram_value[2]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(oram_value[3]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(oram_value[4]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(oram_value[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(oram_value[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(oram_value[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(oram_value[8]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(oram_value[9]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(wb_rst_i),
    .X(net12));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(oram_addr[0]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(oram_addr[1]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(oram_addr[2]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(oram_addr[3]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(oram_addr[4]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(oram_addr[5]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(oram_addr[6]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(oram_addr[7]));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_26 (.LO(net26));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__296__A_N (.DIODE(_045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__254__A (.DIODE(_045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__227__A (.DIODE(_045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__223__A (.DIODE(_045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__219__A (.DIODE(_045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__A (.DIODE(_045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__205__A (.DIODE(_045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A (.DIODE(_045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__166__A (.DIODE(_045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A (.DIODE(_045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__270__A (.DIODE(_054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__267__A (.DIODE(_054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A (.DIODE(_054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__A (.DIODE(_054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__A (.DIODE(_054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__176__A2 (.DIODE(_054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__174__A2 (.DIODE(_054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A1 (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__S1 (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__S1 (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__189__B_N (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__187__A (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__S1 (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__B_N (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__179__A (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__175__S1 (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__173__S1 (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__174__B2 (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__176__B2 (.DIODE(_059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__179__B (.DIODE(_061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__187__B (.DIODE(_063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A (.DIODE(_063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__186__A2 (.DIODE(_066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__189__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A1 (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__196__B2 (.DIODE(_074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__198__B2 (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(oram_value[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(oram_value[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(oram_value[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(oram_value[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(oram_value[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(oram_value[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(oram_value[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(oram_value[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(oram_value[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(oram_value[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(oram_value[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__300__A0 (.DIODE(\tms1x00.PA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__291__A0 (.DIODE(\tms1x00.PA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__229__A1 (.DIODE(\tms1x00.PA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__273__A0 (.DIODE(\tms1x00.PC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__248__A (.DIODE(\tms1x00.PC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__A0 (.DIODE(\tms1x00.PC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__281__A0 (.DIODE(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__266__A1 (.DIODE(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__A0 (.DIODE(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__283__A0 (.DIODE(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__269__A1 (.DIODE(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__A0 (.DIODE(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__234__B_N (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__216__C (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__209__D (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__206__C (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__201__D (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__174__A1 (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__233__A (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__216__B (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__209__C (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__208__A (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__201__C (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__176__A1 (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__293__A (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__262__A1 (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__222__A0 (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__210__C (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__203__A (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A0 (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__294__A (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__A1 (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__226__A0 (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__210__B (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__202__A (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__196__A1 (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__A0 (.DIODE(\tms1x00.ins_in[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__A1 (.DIODE(\tms1x00.ins_in[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__230__A0 (.DIODE(\tms1x00.ins_in[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__210__A (.DIODE(\tms1x00.ins_in[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__204__A0 (.DIODE(\tms1x00.ins_in[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__198__A1 (.DIODE(\tms1x00.ins_in[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__273__A1 (.DIODE(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__S0 (.DIODE(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__S0 (.DIODE(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__S0 (.DIODE(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__188__S (.DIODE(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__S0 (.DIODE(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__180__S (.DIODE(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__178__S (.DIODE(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__175__S0 (.DIODE(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__173__S0 (.DIODE(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__S1 (.DIODE(\tms1x00.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__172__A (.DIODE(\tms1x00.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(wb_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__A3 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__180__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__188__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__188__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__A3 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__A3 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__271__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__C (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__168__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__161__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__156__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_output13_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__199__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_output14_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__206__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__165__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__162__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__160__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_output15_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__271__C (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__206__A_N (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__162__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__160__A_N (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_output16_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__271__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__206__D (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__200__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__170__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__167__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__165__S (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__160__C (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_output17_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_output18_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__277__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_output19_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__279__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_output20_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__281__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__283__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__285__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output23_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__287__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_output24_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__289__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_output25_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__291__A1 (.DIODE(net25));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1378 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1419 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1450 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1480 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1490 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1518 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1524 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1528 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1553 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1574 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1594 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1603 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1618 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1637 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1648 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1659 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1663 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1679 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1689 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1693 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1701 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1706 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1709 ();
 assign io_oeb[0] = net92;
 assign io_oeb[10] = net31;
 assign io_oeb[11] = net32;
 assign io_oeb[12] = net33;
 assign io_oeb[13] = net34;
 assign io_oeb[14] = net35;
 assign io_oeb[15] = net36;
 assign io_oeb[16] = net37;
 assign io_oeb[17] = net38;
 assign io_oeb[18] = net39;
 assign io_oeb[19] = net40;
 assign io_oeb[1] = net93;
 assign io_oeb[20] = net41;
 assign io_oeb[21] = net42;
 assign io_oeb[22] = net43;
 assign io_oeb[23] = net44;
 assign io_oeb[24] = net45;
 assign io_oeb[25] = net46;
 assign io_oeb[26] = net47;
 assign io_oeb[27] = net48;
 assign io_oeb[28] = net49;
 assign io_oeb[29] = net50;
 assign io_oeb[2] = net94;
 assign io_oeb[30] = net51;
 assign io_oeb[31] = net52;
 assign io_oeb[32] = net53;
 assign io_oeb[33] = net54;
 assign io_oeb[34] = net55;
 assign io_oeb[35] = net56;
 assign io_oeb[36] = net57;
 assign io_oeb[37] = net97;
 assign io_oeb[3] = net95;
 assign io_oeb[4] = net96;
 assign io_oeb[5] = net26;
 assign io_oeb[6] = net27;
 assign io_oeb[7] = net28;
 assign io_oeb[8] = net29;
 assign io_oeb[9] = net30;
 assign io_out[0] = net58;
 assign io_out[10] = net68;
 assign io_out[11] = net69;
 assign io_out[12] = net70;
 assign io_out[13] = net71;
 assign io_out[19] = net72;
 assign io_out[1] = net59;
 assign io_out[20] = net73;
 assign io_out[21] = net74;
 assign io_out[22] = net75;
 assign io_out[23] = net76;
 assign io_out[24] = net77;
 assign io_out[25] = net78;
 assign io_out[26] = net79;
 assign io_out[27] = net80;
 assign io_out[28] = net81;
 assign io_out[29] = net82;
 assign io_out[2] = net60;
 assign io_out[30] = net83;
 assign io_out[31] = net84;
 assign io_out[32] = net85;
 assign io_out[33] = net86;
 assign io_out[34] = net87;
 assign io_out[35] = net88;
 assign io_out[36] = net89;
 assign io_out[37] = net90;
 assign io_out[3] = net61;
 assign io_out[4] = net62;
 assign io_out[5] = net63;
 assign io_out[6] = net64;
 assign io_out[7] = net65;
 assign io_out[8] = net66;
 assign io_out[9] = net67;
 assign oram_addr[8] = net91;
endmodule

