magic
tech sky130B
magscale 1 2
timestamp 1679053754
<< obsli1 >>
rect 1104 2159 128892 87601
<< obsm1 >>
rect 934 76 129062 87632
<< metal2 >>
rect 2594 89200 2650 90000
rect 3698 89200 3754 90000
rect 4802 89200 4858 90000
rect 5906 89200 5962 90000
rect 7010 89200 7066 90000
rect 8114 89200 8170 90000
rect 9218 89200 9274 90000
rect 10322 89200 10378 90000
rect 11426 89200 11482 90000
rect 12530 89200 12586 90000
rect 13634 89200 13690 90000
rect 14738 89200 14794 90000
rect 15842 89200 15898 90000
rect 16946 89200 17002 90000
rect 18050 89200 18106 90000
rect 19154 89200 19210 90000
rect 20258 89200 20314 90000
rect 21362 89200 21418 90000
rect 22466 89200 22522 90000
rect 23570 89200 23626 90000
rect 24674 89200 24730 90000
rect 25778 89200 25834 90000
rect 26882 89200 26938 90000
rect 27986 89200 28042 90000
rect 29090 89200 29146 90000
rect 30194 89200 30250 90000
rect 31298 89200 31354 90000
rect 32402 89200 32458 90000
rect 33506 89200 33562 90000
rect 34610 89200 34666 90000
rect 35714 89200 35770 90000
rect 36818 89200 36874 90000
rect 37922 89200 37978 90000
rect 39026 89200 39082 90000
rect 40130 89200 40186 90000
rect 41234 89200 41290 90000
rect 42338 89200 42394 90000
rect 43442 89200 43498 90000
rect 44546 89200 44602 90000
rect 45650 89200 45706 90000
rect 46754 89200 46810 90000
rect 47858 89200 47914 90000
rect 48962 89200 49018 90000
rect 50066 89200 50122 90000
rect 51170 89200 51226 90000
rect 52274 89200 52330 90000
rect 53378 89200 53434 90000
rect 54482 89200 54538 90000
rect 55586 89200 55642 90000
rect 56690 89200 56746 90000
rect 57794 89200 57850 90000
rect 58898 89200 58954 90000
rect 60002 89200 60058 90000
rect 61106 89200 61162 90000
rect 62210 89200 62266 90000
rect 63314 89200 63370 90000
rect 64418 89200 64474 90000
rect 65522 89200 65578 90000
rect 66626 89200 66682 90000
rect 67730 89200 67786 90000
rect 68834 89200 68890 90000
rect 69938 89200 69994 90000
rect 71042 89200 71098 90000
rect 72146 89200 72202 90000
rect 73250 89200 73306 90000
rect 74354 89200 74410 90000
rect 75458 89200 75514 90000
rect 76562 89200 76618 90000
rect 77666 89200 77722 90000
rect 78770 89200 78826 90000
rect 79874 89200 79930 90000
rect 80978 89200 81034 90000
rect 82082 89200 82138 90000
rect 83186 89200 83242 90000
rect 84290 89200 84346 90000
rect 85394 89200 85450 90000
rect 86498 89200 86554 90000
rect 87602 89200 87658 90000
rect 88706 89200 88762 90000
rect 89810 89200 89866 90000
rect 90914 89200 90970 90000
rect 92018 89200 92074 90000
rect 93122 89200 93178 90000
rect 94226 89200 94282 90000
rect 95330 89200 95386 90000
rect 96434 89200 96490 90000
rect 97538 89200 97594 90000
rect 98642 89200 98698 90000
rect 99746 89200 99802 90000
rect 100850 89200 100906 90000
rect 101954 89200 102010 90000
rect 103058 89200 103114 90000
rect 104162 89200 104218 90000
rect 105266 89200 105322 90000
rect 106370 89200 106426 90000
rect 107474 89200 107530 90000
rect 108578 89200 108634 90000
rect 109682 89200 109738 90000
rect 110786 89200 110842 90000
rect 111890 89200 111946 90000
rect 112994 89200 113050 90000
rect 114098 89200 114154 90000
rect 115202 89200 115258 90000
rect 116306 89200 116362 90000
rect 117410 89200 117466 90000
rect 118514 89200 118570 90000
rect 119618 89200 119674 90000
rect 120722 89200 120778 90000
rect 121826 89200 121882 90000
rect 122930 89200 122986 90000
rect 124034 89200 124090 90000
rect 125138 89200 125194 90000
rect 126242 89200 126298 90000
rect 127346 89200 127402 90000
rect 4066 0 4122 800
rect 4894 0 4950 800
rect 5722 0 5778 800
rect 6550 0 6606 800
rect 7378 0 7434 800
rect 8206 0 8262 800
rect 9034 0 9090 800
rect 9862 0 9918 800
rect 10690 0 10746 800
rect 11518 0 11574 800
rect 12346 0 12402 800
rect 13174 0 13230 800
rect 14002 0 14058 800
rect 14830 0 14886 800
rect 15658 0 15714 800
rect 16486 0 16542 800
rect 17314 0 17370 800
rect 18142 0 18198 800
rect 18970 0 19026 800
rect 19798 0 19854 800
rect 20626 0 20682 800
rect 21454 0 21510 800
rect 22282 0 22338 800
rect 23110 0 23166 800
rect 23938 0 23994 800
rect 24766 0 24822 800
rect 25594 0 25650 800
rect 26422 0 26478 800
rect 27250 0 27306 800
rect 28078 0 28134 800
rect 28906 0 28962 800
rect 29734 0 29790 800
rect 30562 0 30618 800
rect 31390 0 31446 800
rect 32218 0 32274 800
rect 33046 0 33102 800
rect 33874 0 33930 800
rect 34702 0 34758 800
rect 35530 0 35586 800
rect 36358 0 36414 800
rect 37186 0 37242 800
rect 38014 0 38070 800
rect 38842 0 38898 800
rect 39670 0 39726 800
rect 40498 0 40554 800
rect 41326 0 41382 800
rect 42154 0 42210 800
rect 42982 0 43038 800
rect 43810 0 43866 800
rect 44638 0 44694 800
rect 45466 0 45522 800
rect 46294 0 46350 800
rect 47122 0 47178 800
rect 47950 0 48006 800
rect 48778 0 48834 800
rect 49606 0 49662 800
rect 50434 0 50490 800
rect 51262 0 51318 800
rect 52090 0 52146 800
rect 52918 0 52974 800
rect 53746 0 53802 800
rect 54574 0 54630 800
rect 55402 0 55458 800
rect 56230 0 56286 800
rect 57058 0 57114 800
rect 57886 0 57942 800
rect 58714 0 58770 800
rect 59542 0 59598 800
rect 60370 0 60426 800
rect 61198 0 61254 800
rect 62026 0 62082 800
rect 62854 0 62910 800
rect 63682 0 63738 800
rect 64510 0 64566 800
rect 65338 0 65394 800
rect 66166 0 66222 800
rect 66994 0 67050 800
rect 67822 0 67878 800
rect 68650 0 68706 800
rect 69478 0 69534 800
rect 70306 0 70362 800
rect 71134 0 71190 800
rect 71962 0 72018 800
rect 72790 0 72846 800
rect 73618 0 73674 800
rect 74446 0 74502 800
rect 75274 0 75330 800
rect 76102 0 76158 800
rect 76930 0 76986 800
rect 77758 0 77814 800
rect 78586 0 78642 800
rect 79414 0 79470 800
rect 80242 0 80298 800
rect 81070 0 81126 800
rect 81898 0 81954 800
rect 82726 0 82782 800
rect 83554 0 83610 800
rect 84382 0 84438 800
rect 85210 0 85266 800
rect 86038 0 86094 800
rect 86866 0 86922 800
rect 87694 0 87750 800
rect 88522 0 88578 800
rect 89350 0 89406 800
rect 90178 0 90234 800
rect 91006 0 91062 800
rect 91834 0 91890 800
rect 92662 0 92718 800
rect 93490 0 93546 800
rect 94318 0 94374 800
rect 95146 0 95202 800
rect 95974 0 96030 800
rect 96802 0 96858 800
rect 97630 0 97686 800
rect 98458 0 98514 800
rect 99286 0 99342 800
rect 100114 0 100170 800
rect 100942 0 100998 800
rect 101770 0 101826 800
rect 102598 0 102654 800
rect 103426 0 103482 800
rect 104254 0 104310 800
rect 105082 0 105138 800
rect 105910 0 105966 800
rect 106738 0 106794 800
rect 107566 0 107622 800
rect 108394 0 108450 800
rect 109222 0 109278 800
rect 110050 0 110106 800
rect 110878 0 110934 800
rect 111706 0 111762 800
rect 112534 0 112590 800
rect 113362 0 113418 800
rect 114190 0 114246 800
rect 115018 0 115074 800
rect 115846 0 115902 800
rect 116674 0 116730 800
rect 117502 0 117558 800
rect 118330 0 118386 800
rect 119158 0 119214 800
rect 119986 0 120042 800
rect 120814 0 120870 800
rect 121642 0 121698 800
rect 122470 0 122526 800
rect 123298 0 123354 800
rect 124126 0 124182 800
rect 124954 0 125010 800
rect 125782 0 125838 800
<< obsm2 >>
rect 938 89144 2538 89298
rect 2706 89144 3642 89298
rect 3810 89144 4746 89298
rect 4914 89144 5850 89298
rect 6018 89144 6954 89298
rect 7122 89144 8058 89298
rect 8226 89144 9162 89298
rect 9330 89144 10266 89298
rect 10434 89144 11370 89298
rect 11538 89144 12474 89298
rect 12642 89144 13578 89298
rect 13746 89144 14682 89298
rect 14850 89144 15786 89298
rect 15954 89144 16890 89298
rect 17058 89144 17994 89298
rect 18162 89144 19098 89298
rect 19266 89144 20202 89298
rect 20370 89144 21306 89298
rect 21474 89144 22410 89298
rect 22578 89144 23514 89298
rect 23682 89144 24618 89298
rect 24786 89144 25722 89298
rect 25890 89144 26826 89298
rect 26994 89144 27930 89298
rect 28098 89144 29034 89298
rect 29202 89144 30138 89298
rect 30306 89144 31242 89298
rect 31410 89144 32346 89298
rect 32514 89144 33450 89298
rect 33618 89144 34554 89298
rect 34722 89144 35658 89298
rect 35826 89144 36762 89298
rect 36930 89144 37866 89298
rect 38034 89144 38970 89298
rect 39138 89144 40074 89298
rect 40242 89144 41178 89298
rect 41346 89144 42282 89298
rect 42450 89144 43386 89298
rect 43554 89144 44490 89298
rect 44658 89144 45594 89298
rect 45762 89144 46698 89298
rect 46866 89144 47802 89298
rect 47970 89144 48906 89298
rect 49074 89144 50010 89298
rect 50178 89144 51114 89298
rect 51282 89144 52218 89298
rect 52386 89144 53322 89298
rect 53490 89144 54426 89298
rect 54594 89144 55530 89298
rect 55698 89144 56634 89298
rect 56802 89144 57738 89298
rect 57906 89144 58842 89298
rect 59010 89144 59946 89298
rect 60114 89144 61050 89298
rect 61218 89144 62154 89298
rect 62322 89144 63258 89298
rect 63426 89144 64362 89298
rect 64530 89144 65466 89298
rect 65634 89144 66570 89298
rect 66738 89144 67674 89298
rect 67842 89144 68778 89298
rect 68946 89144 69882 89298
rect 70050 89144 70986 89298
rect 71154 89144 72090 89298
rect 72258 89144 73194 89298
rect 73362 89144 74298 89298
rect 74466 89144 75402 89298
rect 75570 89144 76506 89298
rect 76674 89144 77610 89298
rect 77778 89144 78714 89298
rect 78882 89144 79818 89298
rect 79986 89144 80922 89298
rect 81090 89144 82026 89298
rect 82194 89144 83130 89298
rect 83298 89144 84234 89298
rect 84402 89144 85338 89298
rect 85506 89144 86442 89298
rect 86610 89144 87546 89298
rect 87714 89144 88650 89298
rect 88818 89144 89754 89298
rect 89922 89144 90858 89298
rect 91026 89144 91962 89298
rect 92130 89144 93066 89298
rect 93234 89144 94170 89298
rect 94338 89144 95274 89298
rect 95442 89144 96378 89298
rect 96546 89144 97482 89298
rect 97650 89144 98586 89298
rect 98754 89144 99690 89298
rect 99858 89144 100794 89298
rect 100962 89144 101898 89298
rect 102066 89144 103002 89298
rect 103170 89144 104106 89298
rect 104274 89144 105210 89298
rect 105378 89144 106314 89298
rect 106482 89144 107418 89298
rect 107586 89144 108522 89298
rect 108690 89144 109626 89298
rect 109794 89144 110730 89298
rect 110898 89144 111834 89298
rect 112002 89144 112938 89298
rect 113106 89144 114042 89298
rect 114210 89144 115146 89298
rect 115314 89144 116250 89298
rect 116418 89144 117354 89298
rect 117522 89144 118458 89298
rect 118626 89144 119562 89298
rect 119730 89144 120666 89298
rect 120834 89144 121770 89298
rect 121938 89144 122874 89298
rect 123042 89144 123978 89298
rect 124146 89144 125082 89298
rect 125250 89144 126186 89298
rect 126354 89144 127290 89298
rect 127458 89144 129058 89298
rect 938 856 129058 89144
rect 938 70 4010 856
rect 4178 70 4838 856
rect 5006 70 5666 856
rect 5834 70 6494 856
rect 6662 70 7322 856
rect 7490 70 8150 856
rect 8318 70 8978 856
rect 9146 70 9806 856
rect 9974 70 10634 856
rect 10802 70 11462 856
rect 11630 70 12290 856
rect 12458 70 13118 856
rect 13286 70 13946 856
rect 14114 70 14774 856
rect 14942 70 15602 856
rect 15770 70 16430 856
rect 16598 70 17258 856
rect 17426 70 18086 856
rect 18254 70 18914 856
rect 19082 70 19742 856
rect 19910 70 20570 856
rect 20738 70 21398 856
rect 21566 70 22226 856
rect 22394 70 23054 856
rect 23222 70 23882 856
rect 24050 70 24710 856
rect 24878 70 25538 856
rect 25706 70 26366 856
rect 26534 70 27194 856
rect 27362 70 28022 856
rect 28190 70 28850 856
rect 29018 70 29678 856
rect 29846 70 30506 856
rect 30674 70 31334 856
rect 31502 70 32162 856
rect 32330 70 32990 856
rect 33158 70 33818 856
rect 33986 70 34646 856
rect 34814 70 35474 856
rect 35642 70 36302 856
rect 36470 70 37130 856
rect 37298 70 37958 856
rect 38126 70 38786 856
rect 38954 70 39614 856
rect 39782 70 40442 856
rect 40610 70 41270 856
rect 41438 70 42098 856
rect 42266 70 42926 856
rect 43094 70 43754 856
rect 43922 70 44582 856
rect 44750 70 45410 856
rect 45578 70 46238 856
rect 46406 70 47066 856
rect 47234 70 47894 856
rect 48062 70 48722 856
rect 48890 70 49550 856
rect 49718 70 50378 856
rect 50546 70 51206 856
rect 51374 70 52034 856
rect 52202 70 52862 856
rect 53030 70 53690 856
rect 53858 70 54518 856
rect 54686 70 55346 856
rect 55514 70 56174 856
rect 56342 70 57002 856
rect 57170 70 57830 856
rect 57998 70 58658 856
rect 58826 70 59486 856
rect 59654 70 60314 856
rect 60482 70 61142 856
rect 61310 70 61970 856
rect 62138 70 62798 856
rect 62966 70 63626 856
rect 63794 70 64454 856
rect 64622 70 65282 856
rect 65450 70 66110 856
rect 66278 70 66938 856
rect 67106 70 67766 856
rect 67934 70 68594 856
rect 68762 70 69422 856
rect 69590 70 70250 856
rect 70418 70 71078 856
rect 71246 70 71906 856
rect 72074 70 72734 856
rect 72902 70 73562 856
rect 73730 70 74390 856
rect 74558 70 75218 856
rect 75386 70 76046 856
rect 76214 70 76874 856
rect 77042 70 77702 856
rect 77870 70 78530 856
rect 78698 70 79358 856
rect 79526 70 80186 856
rect 80354 70 81014 856
rect 81182 70 81842 856
rect 82010 70 82670 856
rect 82838 70 83498 856
rect 83666 70 84326 856
rect 84494 70 85154 856
rect 85322 70 85982 856
rect 86150 70 86810 856
rect 86978 70 87638 856
rect 87806 70 88466 856
rect 88634 70 89294 856
rect 89462 70 90122 856
rect 90290 70 90950 856
rect 91118 70 91778 856
rect 91946 70 92606 856
rect 92774 70 93434 856
rect 93602 70 94262 856
rect 94430 70 95090 856
rect 95258 70 95918 856
rect 96086 70 96746 856
rect 96914 70 97574 856
rect 97742 70 98402 856
rect 98570 70 99230 856
rect 99398 70 100058 856
rect 100226 70 100886 856
rect 101054 70 101714 856
rect 101882 70 102542 856
rect 102710 70 103370 856
rect 103538 70 104198 856
rect 104366 70 105026 856
rect 105194 70 105854 856
rect 106022 70 106682 856
rect 106850 70 107510 856
rect 107678 70 108338 856
rect 108506 70 109166 856
rect 109334 70 109994 856
rect 110162 70 110822 856
rect 110990 70 111650 856
rect 111818 70 112478 856
rect 112646 70 113306 856
rect 113474 70 114134 856
rect 114302 70 114962 856
rect 115130 70 115790 856
rect 115958 70 116618 856
rect 116786 70 117446 856
rect 117614 70 118274 856
rect 118442 70 119102 856
rect 119270 70 119930 856
rect 120098 70 120758 856
rect 120926 70 121586 856
rect 121754 70 122414 856
rect 122582 70 123242 856
rect 123410 70 124070 856
rect 124238 70 124898 856
rect 125066 70 125726 856
rect 125894 70 129058 856
<< metal3 >>
rect 0 86776 800 86896
rect 129200 86776 130000 86896
rect 0 84736 800 84856
rect 0 82696 800 82816
rect 129200 81200 130000 81320
rect 0 80656 800 80776
rect 0 78616 800 78736
rect 0 76576 800 76696
rect 129200 75624 130000 75744
rect 0 74536 800 74656
rect 0 72496 800 72616
rect 0 70456 800 70576
rect 129200 70048 130000 70168
rect 0 68416 800 68536
rect 0 66376 800 66496
rect 0 64336 800 64456
rect 129200 64472 130000 64592
rect 0 62296 800 62416
rect 0 60256 800 60376
rect 129200 58896 130000 59016
rect 0 58216 800 58336
rect 0 56176 800 56296
rect 0 54136 800 54256
rect 129200 53320 130000 53440
rect 0 52096 800 52216
rect 0 50056 800 50176
rect 0 48016 800 48136
rect 129200 47744 130000 47864
rect 0 45976 800 46096
rect 0 43936 800 44056
rect 129200 42168 130000 42288
rect 0 41896 800 42016
rect 0 39856 800 39976
rect 0 37816 800 37936
rect 129200 36592 130000 36712
rect 0 35776 800 35896
rect 0 33736 800 33856
rect 0 31696 800 31816
rect 129200 31016 130000 31136
rect 0 29656 800 29776
rect 0 27616 800 27736
rect 0 25576 800 25696
rect 129200 25440 130000 25560
rect 0 23536 800 23656
rect 0 21496 800 21616
rect 129200 19864 130000 19984
rect 0 19456 800 19576
rect 0 17416 800 17536
rect 0 15376 800 15496
rect 129200 14288 130000 14408
rect 0 13336 800 13456
rect 0 11296 800 11416
rect 0 9256 800 9376
rect 129200 8712 130000 8832
rect 0 7216 800 7336
rect 0 5176 800 5296
rect 0 3136 800 3256
rect 129200 3136 130000 3256
<< obsm3 >>
rect 800 86976 129200 87617
rect 880 86696 129120 86976
rect 800 84936 129200 86696
rect 880 84656 129200 84936
rect 800 82896 129200 84656
rect 880 82616 129200 82896
rect 800 81400 129200 82616
rect 800 81120 129120 81400
rect 800 80856 129200 81120
rect 880 80576 129200 80856
rect 800 78816 129200 80576
rect 880 78536 129200 78816
rect 800 76776 129200 78536
rect 880 76496 129200 76776
rect 800 75824 129200 76496
rect 800 75544 129120 75824
rect 800 74736 129200 75544
rect 880 74456 129200 74736
rect 800 72696 129200 74456
rect 880 72416 129200 72696
rect 800 70656 129200 72416
rect 880 70376 129200 70656
rect 800 70248 129200 70376
rect 800 69968 129120 70248
rect 800 68616 129200 69968
rect 880 68336 129200 68616
rect 800 66576 129200 68336
rect 880 66296 129200 66576
rect 800 64672 129200 66296
rect 800 64536 129120 64672
rect 880 64392 129120 64536
rect 880 64256 129200 64392
rect 800 62496 129200 64256
rect 880 62216 129200 62496
rect 800 60456 129200 62216
rect 880 60176 129200 60456
rect 800 59096 129200 60176
rect 800 58816 129120 59096
rect 800 58416 129200 58816
rect 880 58136 129200 58416
rect 800 56376 129200 58136
rect 880 56096 129200 56376
rect 800 54336 129200 56096
rect 880 54056 129200 54336
rect 800 53520 129200 54056
rect 800 53240 129120 53520
rect 800 52296 129200 53240
rect 880 52016 129200 52296
rect 800 50256 129200 52016
rect 880 49976 129200 50256
rect 800 48216 129200 49976
rect 880 47944 129200 48216
rect 880 47936 129120 47944
rect 800 47664 129120 47936
rect 800 46176 129200 47664
rect 880 45896 129200 46176
rect 800 44136 129200 45896
rect 880 43856 129200 44136
rect 800 42368 129200 43856
rect 800 42096 129120 42368
rect 880 42088 129120 42096
rect 880 41816 129200 42088
rect 800 40056 129200 41816
rect 880 39776 129200 40056
rect 800 38016 129200 39776
rect 880 37736 129200 38016
rect 800 36792 129200 37736
rect 800 36512 129120 36792
rect 800 35976 129200 36512
rect 880 35696 129200 35976
rect 800 33936 129200 35696
rect 880 33656 129200 33936
rect 800 31896 129200 33656
rect 880 31616 129200 31896
rect 800 31216 129200 31616
rect 800 30936 129120 31216
rect 800 29856 129200 30936
rect 880 29576 129200 29856
rect 800 27816 129200 29576
rect 880 27536 129200 27816
rect 800 25776 129200 27536
rect 880 25640 129200 25776
rect 880 25496 129120 25640
rect 800 25360 129120 25496
rect 800 23736 129200 25360
rect 880 23456 129200 23736
rect 800 21696 129200 23456
rect 880 21416 129200 21696
rect 800 20064 129200 21416
rect 800 19784 129120 20064
rect 800 19656 129200 19784
rect 880 19376 129200 19656
rect 800 17616 129200 19376
rect 880 17336 129200 17616
rect 800 15576 129200 17336
rect 880 15296 129200 15576
rect 800 14488 129200 15296
rect 800 14208 129120 14488
rect 800 13536 129200 14208
rect 880 13256 129200 13536
rect 800 11496 129200 13256
rect 880 11216 129200 11496
rect 800 9456 129200 11216
rect 880 9176 129200 9456
rect 800 8912 129200 9176
rect 800 8632 129120 8912
rect 800 7416 129200 8632
rect 880 7136 129200 7416
rect 800 5376 129200 7136
rect 880 5096 129200 5376
rect 800 3336 129200 5096
rect 880 3056 129120 3336
rect 800 1667 129200 3056
<< metal4 >>
rect 4208 2128 4528 87632
rect 19568 2128 19888 87632
rect 34928 2128 35248 87632
rect 50288 2128 50608 87632
rect 65648 2128 65968 87632
rect 81008 2128 81328 87632
rect 96368 2128 96688 87632
rect 111728 2128 112048 87632
rect 127088 2128 127408 87632
<< obsm4 >>
rect 1899 2619 4128 87413
rect 4608 2619 19488 87413
rect 19968 2619 34848 87413
rect 35328 2619 50208 87413
rect 50688 2619 65568 87413
rect 66048 2619 80928 87413
rect 81408 2619 96288 87413
rect 96768 2619 111648 87413
rect 112128 2619 117885 87413
<< labels >>
rlabel metal2 s 2594 89200 2650 90000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 35714 89200 35770 90000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 39026 89200 39082 90000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 42338 89200 42394 90000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 45650 89200 45706 90000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 48962 89200 49018 90000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 52274 89200 52330 90000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 55586 89200 55642 90000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 58898 89200 58954 90000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 62210 89200 62266 90000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 65522 89200 65578 90000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5906 89200 5962 90000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 68834 89200 68890 90000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 72146 89200 72202 90000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 75458 89200 75514 90000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 78770 89200 78826 90000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 82082 89200 82138 90000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 85394 89200 85450 90000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 88706 89200 88762 90000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 92018 89200 92074 90000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 95330 89200 95386 90000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 98642 89200 98698 90000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 9218 89200 9274 90000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 101954 89200 102010 90000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 105266 89200 105322 90000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 108578 89200 108634 90000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 111890 89200 111946 90000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 115202 89200 115258 90000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 118514 89200 118570 90000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 121826 89200 121882 90000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 125138 89200 125194 90000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 12530 89200 12586 90000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 15842 89200 15898 90000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 19154 89200 19210 90000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 22466 89200 22522 90000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 25778 89200 25834 90000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 29090 89200 29146 90000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 32402 89200 32458 90000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3698 89200 3754 90000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 36818 89200 36874 90000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 40130 89200 40186 90000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 43442 89200 43498 90000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 46754 89200 46810 90000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 50066 89200 50122 90000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 53378 89200 53434 90000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 56690 89200 56746 90000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 60002 89200 60058 90000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 63314 89200 63370 90000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 66626 89200 66682 90000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7010 89200 7066 90000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 69938 89200 69994 90000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 73250 89200 73306 90000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 76562 89200 76618 90000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 79874 89200 79930 90000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 83186 89200 83242 90000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 86498 89200 86554 90000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 89810 89200 89866 90000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 93122 89200 93178 90000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 96434 89200 96490 90000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 99746 89200 99802 90000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 10322 89200 10378 90000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 103058 89200 103114 90000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 106370 89200 106426 90000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 109682 89200 109738 90000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 112994 89200 113050 90000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 116306 89200 116362 90000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 119618 89200 119674 90000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 122930 89200 122986 90000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 126242 89200 126298 90000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 13634 89200 13690 90000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 16946 89200 17002 90000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 20258 89200 20314 90000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 23570 89200 23626 90000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 26882 89200 26938 90000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 30194 89200 30250 90000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 33506 89200 33562 90000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4802 89200 4858 90000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 37922 89200 37978 90000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 41234 89200 41290 90000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 44546 89200 44602 90000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 47858 89200 47914 90000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 51170 89200 51226 90000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 54482 89200 54538 90000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 57794 89200 57850 90000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 61106 89200 61162 90000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 64418 89200 64474 90000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 67730 89200 67786 90000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8114 89200 8170 90000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 71042 89200 71098 90000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 74354 89200 74410 90000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 77666 89200 77722 90000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 80978 89200 81034 90000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 84290 89200 84346 90000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 87602 89200 87658 90000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 90914 89200 90970 90000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 94226 89200 94282 90000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 97538 89200 97594 90000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 100850 89200 100906 90000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 11426 89200 11482 90000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 104162 89200 104218 90000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 107474 89200 107530 90000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 110786 89200 110842 90000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 114098 89200 114154 90000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 117410 89200 117466 90000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 120722 89200 120778 90000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 124034 89200 124090 90000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 127346 89200 127402 90000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 14738 89200 14794 90000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 18050 89200 18106 90000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 21362 89200 21418 90000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 24674 89200 24730 90000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 27986 89200 28042 90000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 31298 89200 31354 90000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 34610 89200 34666 90000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 129200 8712 130000 8832 6 ram_addr[0]
port 118 nsew signal output
rlabel metal3 s 129200 25440 130000 25560 6 ram_addr[1]
port 119 nsew signal output
rlabel metal3 s 129200 42168 130000 42288 6 ram_addr[2]
port 120 nsew signal output
rlabel metal3 s 129200 58896 130000 59016 6 ram_addr[3]
port 121 nsew signal output
rlabel metal3 s 129200 75624 130000 75744 6 ram_addr[4]
port 122 nsew signal output
rlabel metal3 s 129200 81200 130000 81320 6 ram_addr[5]
port 123 nsew signal output
rlabel metal3 s 129200 86776 130000 86896 6 ram_addr[6]
port 124 nsew signal output
rlabel metal3 s 129200 14288 130000 14408 6 ram_val_in[0]
port 125 nsew signal input
rlabel metal3 s 129200 31016 130000 31136 6 ram_val_in[1]
port 126 nsew signal input
rlabel metal3 s 129200 47744 130000 47864 6 ram_val_in[2]
port 127 nsew signal input
rlabel metal3 s 129200 64472 130000 64592 6 ram_val_in[3]
port 128 nsew signal input
rlabel metal3 s 129200 19864 130000 19984 6 ram_val_out[0]
port 129 nsew signal output
rlabel metal3 s 129200 36592 130000 36712 6 ram_val_out[1]
port 130 nsew signal output
rlabel metal3 s 129200 53320 130000 53440 6 ram_val_out[2]
port 131 nsew signal output
rlabel metal3 s 129200 70048 130000 70168 6 ram_val_out[3]
port 132 nsew signal output
rlabel metal3 s 129200 3136 130000 3256 6 ram_we
port 133 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 rom_addr[0]
port 134 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 rom_addr[1]
port 135 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 rom_addr[2]
port 136 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 rom_addr[3]
port 137 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 rom_addr[4]
port 138 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 rom_addr[5]
port 139 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 rom_addr[6]
port 140 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 rom_addr[7]
port 141 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 rom_addr[8]
port 142 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 rom_csb
port 143 nsew signal output
rlabel metal3 s 0 7216 800 7336 6 rom_value[0]
port 144 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 rom_value[10]
port 145 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 rom_value[11]
port 146 nsew signal input
rlabel metal3 s 0 48016 800 48136 6 rom_value[12]
port 147 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 rom_value[13]
port 148 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 rom_value[14]
port 149 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 rom_value[15]
port 150 nsew signal input
rlabel metal3 s 0 56176 800 56296 6 rom_value[16]
port 151 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 rom_value[17]
port 152 nsew signal input
rlabel metal3 s 0 60256 800 60376 6 rom_value[18]
port 153 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 rom_value[19]
port 154 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 rom_value[1]
port 155 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 rom_value[20]
port 156 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 rom_value[21]
port 157 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 rom_value[22]
port 158 nsew signal input
rlabel metal3 s 0 70456 800 70576 6 rom_value[23]
port 159 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 rom_value[24]
port 160 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 rom_value[25]
port 161 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 rom_value[26]
port 162 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 rom_value[27]
port 163 nsew signal input
rlabel metal3 s 0 80656 800 80776 6 rom_value[28]
port 164 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 rom_value[29]
port 165 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 rom_value[2]
port 166 nsew signal input
rlabel metal3 s 0 84736 800 84856 6 rom_value[30]
port 167 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 rom_value[31]
port 168 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 rom_value[3]
port 169 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 rom_value[4]
port 170 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 rom_value[5]
port 171 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 rom_value[6]
port 172 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 rom_value[7]
port 173 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 rom_value[8]
port 174 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 rom_value[9]
port 175 nsew signal input
rlabel metal4 s 4208 2128 4528 87632 6 vccd1
port 176 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 87632 6 vccd1
port 176 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 87632 6 vccd1
port 176 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 87632 6 vccd1
port 176 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 87632 6 vccd1
port 176 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 87632 6 vssd1
port 177 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 87632 6 vssd1
port 177 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 87632 6 vssd1
port 177 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 87632 6 vssd1
port 177 nsew ground bidirectional
rlabel metal2 s 4066 0 4122 800 6 wb_clk_i
port 178 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wb_rom_adrb[0]
port 179 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wb_rom_adrb[1]
port 180 nsew signal output
rlabel metal2 s 10690 0 10746 800 6 wb_rom_adrb[2]
port 181 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wb_rom_adrb[3]
port 182 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wb_rom_adrb[4]
port 183 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 wb_rom_adrb[5]
port 184 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wb_rom_adrb[6]
port 185 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wb_rom_adrb[7]
port 186 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wb_rom_adrb[8]
port 187 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wb_rom_csb
port 188 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 wb_rom_val[0]
port 189 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wb_rom_val[10]
port 190 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wb_rom_val[11]
port 191 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wb_rom_val[12]
port 192 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wb_rom_val[13]
port 193 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wb_rom_val[14]
port 194 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wb_rom_val[15]
port 195 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wb_rom_val[16]
port 196 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wb_rom_val[17]
port 197 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wb_rom_val[18]
port 198 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wb_rom_val[19]
port 199 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wb_rom_val[1]
port 200 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wb_rom_val[20]
port 201 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wb_rom_val[21]
port 202 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wb_rom_val[22]
port 203 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wb_rom_val[23]
port 204 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wb_rom_val[24]
port 205 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wb_rom_val[25]
port 206 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wb_rom_val[26]
port 207 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wb_rom_val[27]
port 208 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wb_rom_val[28]
port 209 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 wb_rom_val[29]
port 210 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wb_rom_val[2]
port 211 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wb_rom_val[30]
port 212 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wb_rom_val[31]
port 213 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wb_rom_val[3]
port 214 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wb_rom_val[4]
port 215 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wb_rom_val[5]
port 216 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wb_rom_val[6]
port 217 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wb_rom_val[7]
port 218 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wb_rom_val[8]
port 219 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wb_rom_val[9]
port 220 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wb_rom_web
port 221 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wb_rst_i
port 222 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_ack_o
port 223 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 wbs_adr_i[0]
port 224 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 wbs_adr_i[10]
port 225 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 wbs_adr_i[11]
port 226 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 wbs_adr_i[12]
port 227 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 wbs_adr_i[13]
port 228 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 wbs_adr_i[14]
port 229 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 wbs_adr_i[15]
port 230 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 wbs_adr_i[16]
port 231 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 wbs_adr_i[17]
port 232 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 wbs_adr_i[18]
port 233 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 wbs_adr_i[19]
port 234 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_adr_i[1]
port 235 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 wbs_adr_i[20]
port 236 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 wbs_adr_i[21]
port 237 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 wbs_adr_i[22]
port 238 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 wbs_adr_i[23]
port 239 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 wbs_adr_i[24]
port 240 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 wbs_adr_i[25]
port 241 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 wbs_adr_i[26]
port 242 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 wbs_adr_i[27]
port 243 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 wbs_adr_i[28]
port 244 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 wbs_adr_i[29]
port 245 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_adr_i[2]
port 246 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 wbs_adr_i[30]
port 247 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 wbs_adr_i[31]
port 248 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 wbs_adr_i[3]
port 249 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 wbs_adr_i[4]
port 250 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 wbs_adr_i[5]
port 251 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 wbs_adr_i[6]
port 252 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 wbs_adr_i[7]
port 253 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 wbs_adr_i[8]
port 254 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 wbs_adr_i[9]
port 255 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_cyc_i
port 256 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_i[0]
port 257 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 wbs_dat_i[10]
port 258 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 wbs_dat_i[11]
port 259 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 wbs_dat_i[12]
port 260 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 wbs_dat_i[13]
port 261 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 wbs_dat_i[14]
port 262 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 wbs_dat_i[15]
port 263 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 wbs_dat_i[16]
port 264 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 wbs_dat_i[17]
port 265 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 wbs_dat_i[18]
port 266 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 wbs_dat_i[19]
port 267 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 wbs_dat_i[1]
port 268 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 wbs_dat_i[20]
port 269 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 wbs_dat_i[21]
port 270 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 wbs_dat_i[22]
port 271 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 wbs_dat_i[23]
port 272 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 wbs_dat_i[24]
port 273 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 wbs_dat_i[25]
port 274 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 wbs_dat_i[26]
port 275 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 wbs_dat_i[27]
port 276 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 wbs_dat_i[28]
port 277 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 wbs_dat_i[29]
port 278 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_dat_i[2]
port 279 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 wbs_dat_i[30]
port 280 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 wbs_dat_i[31]
port 281 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 wbs_dat_i[3]
port 282 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_dat_i[4]
port 283 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 wbs_dat_i[5]
port 284 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 wbs_dat_i[6]
port 285 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 wbs_dat_i[7]
port 286 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_i[8]
port 287 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 wbs_dat_i[9]
port 288 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 wbs_dat_o[0]
port 289 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 wbs_dat_o[10]
port 290 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 wbs_dat_o[11]
port 291 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 wbs_dat_o[12]
port 292 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 wbs_dat_o[13]
port 293 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 wbs_dat_o[14]
port 294 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 wbs_dat_o[15]
port 295 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 wbs_dat_o[16]
port 296 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 wbs_dat_o[17]
port 297 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 wbs_dat_o[18]
port 298 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 wbs_dat_o[19]
port 299 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 wbs_dat_o[1]
port 300 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 wbs_dat_o[20]
port 301 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 wbs_dat_o[21]
port 302 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 wbs_dat_o[22]
port 303 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 wbs_dat_o[23]
port 304 nsew signal output
rlabel metal2 s 105910 0 105966 800 6 wbs_dat_o[24]
port 305 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 wbs_dat_o[25]
port 306 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 wbs_dat_o[26]
port 307 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 wbs_dat_o[27]
port 308 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 wbs_dat_o[28]
port 309 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 wbs_dat_o[29]
port 310 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_o[2]
port 311 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 wbs_dat_o[30]
port 312 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 wbs_dat_o[31]
port 313 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_o[3]
port 314 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 wbs_dat_o[4]
port 315 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_o[5]
port 316 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 wbs_dat_o[6]
port 317 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 wbs_dat_o[7]
port 318 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 wbs_dat_o[8]
port 319 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 wbs_dat_o[9]
port 320 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_stb_i
port 321 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_we_i
port 322 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 130000 90000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 26346268
string GDS_FILE /home/lucah/mpw-8-as1x00/openlane/wrapped_tms1x00/runs/23_03_17_12_34/results/signoff/wrapped_tms1x00.magic.gds
string GDS_START 967036
<< end >>

