// This is the unpowered netlist.
module wrapped_tms1x00 (oram_csb,
    ram_csb,
    ram_web,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    oram_addr,
    oram_value,
    ram_adrb,
    ram_val,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 output oram_csb;
 output ram_csb;
 output ram_web;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [8:0] oram_addr;
 input [31:0] oram_value;
 output [8:0] ram_adrb;
 input [31:0] ram_val;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire \K_override[0] ;
 wire \K_override[1] ;
 wire \K_override[2] ;
 wire \K_override[3] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire chip_sel_override;
 wire feedback_delay;
 wire net195;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net196;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net197;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire clknet_leaf_0_wb_clk_i;
 wire net182;
 wire net183;
 wire net184;
 wire net192;
 wire net193;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net194;
 wire \tms1x00.A[0] ;
 wire \tms1x00.A[1] ;
 wire \tms1x00.A[2] ;
 wire \tms1x00.A[3] ;
 wire \tms1x00.CL ;
 wire \tms1x00.K_in[0] ;
 wire \tms1x00.K_in[1] ;
 wire \tms1x00.K_in[2] ;
 wire \tms1x00.K_in[3] ;
 wire \tms1x00.K_latch[0] ;
 wire \tms1x00.K_latch[1] ;
 wire \tms1x00.K_latch[2] ;
 wire \tms1x00.K_latch[3] ;
 wire \tms1x00.N[0] ;
 wire \tms1x00.N[1] ;
 wire \tms1x00.N[2] ;
 wire \tms1x00.N[3] ;
 wire \tms1x00.PA[0] ;
 wire \tms1x00.PA[1] ;
 wire \tms1x00.PA[2] ;
 wire \tms1x00.PA[3] ;
 wire \tms1x00.PB[0] ;
 wire \tms1x00.PB[1] ;
 wire \tms1x00.PB[2] ;
 wire \tms1x00.PB[3] ;
 wire \tms1x00.PC[0] ;
 wire \tms1x00.PC[1] ;
 wire \tms1x00.PC[2] ;
 wire \tms1x00.PC[3] ;
 wire \tms1x00.PC[4] ;
 wire \tms1x00.PC[5] ;
 wire \tms1x00.P[0] ;
 wire \tms1x00.P[1] ;
 wire \tms1x00.P[2] ;
 wire \tms1x00.P[3] ;
 wire \tms1x00.RAM[0][0] ;
 wire \tms1x00.RAM[0][1] ;
 wire \tms1x00.RAM[0][2] ;
 wire \tms1x00.RAM[0][3] ;
 wire \tms1x00.RAM[100][0] ;
 wire \tms1x00.RAM[100][1] ;
 wire \tms1x00.RAM[100][2] ;
 wire \tms1x00.RAM[100][3] ;
 wire \tms1x00.RAM[101][0] ;
 wire \tms1x00.RAM[101][1] ;
 wire \tms1x00.RAM[101][2] ;
 wire \tms1x00.RAM[101][3] ;
 wire \tms1x00.RAM[102][0] ;
 wire \tms1x00.RAM[102][1] ;
 wire \tms1x00.RAM[102][2] ;
 wire \tms1x00.RAM[102][3] ;
 wire \tms1x00.RAM[103][0] ;
 wire \tms1x00.RAM[103][1] ;
 wire \tms1x00.RAM[103][2] ;
 wire \tms1x00.RAM[103][3] ;
 wire \tms1x00.RAM[104][0] ;
 wire \tms1x00.RAM[104][1] ;
 wire \tms1x00.RAM[104][2] ;
 wire \tms1x00.RAM[104][3] ;
 wire \tms1x00.RAM[105][0] ;
 wire \tms1x00.RAM[105][1] ;
 wire \tms1x00.RAM[105][2] ;
 wire \tms1x00.RAM[105][3] ;
 wire \tms1x00.RAM[106][0] ;
 wire \tms1x00.RAM[106][1] ;
 wire \tms1x00.RAM[106][2] ;
 wire \tms1x00.RAM[106][3] ;
 wire \tms1x00.RAM[107][0] ;
 wire \tms1x00.RAM[107][1] ;
 wire \tms1x00.RAM[107][2] ;
 wire \tms1x00.RAM[107][3] ;
 wire \tms1x00.RAM[108][0] ;
 wire \tms1x00.RAM[108][1] ;
 wire \tms1x00.RAM[108][2] ;
 wire \tms1x00.RAM[108][3] ;
 wire \tms1x00.RAM[109][0] ;
 wire \tms1x00.RAM[109][1] ;
 wire \tms1x00.RAM[109][2] ;
 wire \tms1x00.RAM[109][3] ;
 wire \tms1x00.RAM[10][0] ;
 wire \tms1x00.RAM[10][1] ;
 wire \tms1x00.RAM[10][2] ;
 wire \tms1x00.RAM[10][3] ;
 wire \tms1x00.RAM[110][0] ;
 wire \tms1x00.RAM[110][1] ;
 wire \tms1x00.RAM[110][2] ;
 wire \tms1x00.RAM[110][3] ;
 wire \tms1x00.RAM[111][0] ;
 wire \tms1x00.RAM[111][1] ;
 wire \tms1x00.RAM[111][2] ;
 wire \tms1x00.RAM[111][3] ;
 wire \tms1x00.RAM[112][0] ;
 wire \tms1x00.RAM[112][1] ;
 wire \tms1x00.RAM[112][2] ;
 wire \tms1x00.RAM[112][3] ;
 wire \tms1x00.RAM[113][0] ;
 wire \tms1x00.RAM[113][1] ;
 wire \tms1x00.RAM[113][2] ;
 wire \tms1x00.RAM[113][3] ;
 wire \tms1x00.RAM[114][0] ;
 wire \tms1x00.RAM[114][1] ;
 wire \tms1x00.RAM[114][2] ;
 wire \tms1x00.RAM[114][3] ;
 wire \tms1x00.RAM[115][0] ;
 wire \tms1x00.RAM[115][1] ;
 wire \tms1x00.RAM[115][2] ;
 wire \tms1x00.RAM[115][3] ;
 wire \tms1x00.RAM[116][0] ;
 wire \tms1x00.RAM[116][1] ;
 wire \tms1x00.RAM[116][2] ;
 wire \tms1x00.RAM[116][3] ;
 wire \tms1x00.RAM[117][0] ;
 wire \tms1x00.RAM[117][1] ;
 wire \tms1x00.RAM[117][2] ;
 wire \tms1x00.RAM[117][3] ;
 wire \tms1x00.RAM[118][0] ;
 wire \tms1x00.RAM[118][1] ;
 wire \tms1x00.RAM[118][2] ;
 wire \tms1x00.RAM[118][3] ;
 wire \tms1x00.RAM[119][0] ;
 wire \tms1x00.RAM[119][1] ;
 wire \tms1x00.RAM[119][2] ;
 wire \tms1x00.RAM[119][3] ;
 wire \tms1x00.RAM[11][0] ;
 wire \tms1x00.RAM[11][1] ;
 wire \tms1x00.RAM[11][2] ;
 wire \tms1x00.RAM[11][3] ;
 wire \tms1x00.RAM[120][0] ;
 wire \tms1x00.RAM[120][1] ;
 wire \tms1x00.RAM[120][2] ;
 wire \tms1x00.RAM[120][3] ;
 wire \tms1x00.RAM[121][0] ;
 wire \tms1x00.RAM[121][1] ;
 wire \tms1x00.RAM[121][2] ;
 wire \tms1x00.RAM[121][3] ;
 wire \tms1x00.RAM[122][0] ;
 wire \tms1x00.RAM[122][1] ;
 wire \tms1x00.RAM[122][2] ;
 wire \tms1x00.RAM[122][3] ;
 wire \tms1x00.RAM[123][0] ;
 wire \tms1x00.RAM[123][1] ;
 wire \tms1x00.RAM[123][2] ;
 wire \tms1x00.RAM[123][3] ;
 wire \tms1x00.RAM[124][0] ;
 wire \tms1x00.RAM[124][1] ;
 wire \tms1x00.RAM[124][2] ;
 wire \tms1x00.RAM[124][3] ;
 wire \tms1x00.RAM[125][0] ;
 wire \tms1x00.RAM[125][1] ;
 wire \tms1x00.RAM[125][2] ;
 wire \tms1x00.RAM[125][3] ;
 wire \tms1x00.RAM[126][0] ;
 wire \tms1x00.RAM[126][1] ;
 wire \tms1x00.RAM[126][2] ;
 wire \tms1x00.RAM[126][3] ;
 wire \tms1x00.RAM[127][0] ;
 wire \tms1x00.RAM[127][1] ;
 wire \tms1x00.RAM[127][2] ;
 wire \tms1x00.RAM[127][3] ;
 wire \tms1x00.RAM[12][0] ;
 wire \tms1x00.RAM[12][1] ;
 wire \tms1x00.RAM[12][2] ;
 wire \tms1x00.RAM[12][3] ;
 wire \tms1x00.RAM[13][0] ;
 wire \tms1x00.RAM[13][1] ;
 wire \tms1x00.RAM[13][2] ;
 wire \tms1x00.RAM[13][3] ;
 wire \tms1x00.RAM[14][0] ;
 wire \tms1x00.RAM[14][1] ;
 wire \tms1x00.RAM[14][2] ;
 wire \tms1x00.RAM[14][3] ;
 wire \tms1x00.RAM[15][0] ;
 wire \tms1x00.RAM[15][1] ;
 wire \tms1x00.RAM[15][2] ;
 wire \tms1x00.RAM[15][3] ;
 wire \tms1x00.RAM[16][0] ;
 wire \tms1x00.RAM[16][1] ;
 wire \tms1x00.RAM[16][2] ;
 wire \tms1x00.RAM[16][3] ;
 wire \tms1x00.RAM[17][0] ;
 wire \tms1x00.RAM[17][1] ;
 wire \tms1x00.RAM[17][2] ;
 wire \tms1x00.RAM[17][3] ;
 wire \tms1x00.RAM[18][0] ;
 wire \tms1x00.RAM[18][1] ;
 wire \tms1x00.RAM[18][2] ;
 wire \tms1x00.RAM[18][3] ;
 wire \tms1x00.RAM[19][0] ;
 wire \tms1x00.RAM[19][1] ;
 wire \tms1x00.RAM[19][2] ;
 wire \tms1x00.RAM[19][3] ;
 wire \tms1x00.RAM[1][0] ;
 wire \tms1x00.RAM[1][1] ;
 wire \tms1x00.RAM[1][2] ;
 wire \tms1x00.RAM[1][3] ;
 wire \tms1x00.RAM[20][0] ;
 wire \tms1x00.RAM[20][1] ;
 wire \tms1x00.RAM[20][2] ;
 wire \tms1x00.RAM[20][3] ;
 wire \tms1x00.RAM[21][0] ;
 wire \tms1x00.RAM[21][1] ;
 wire \tms1x00.RAM[21][2] ;
 wire \tms1x00.RAM[21][3] ;
 wire \tms1x00.RAM[22][0] ;
 wire \tms1x00.RAM[22][1] ;
 wire \tms1x00.RAM[22][2] ;
 wire \tms1x00.RAM[22][3] ;
 wire \tms1x00.RAM[23][0] ;
 wire \tms1x00.RAM[23][1] ;
 wire \tms1x00.RAM[23][2] ;
 wire \tms1x00.RAM[23][3] ;
 wire \tms1x00.RAM[24][0] ;
 wire \tms1x00.RAM[24][1] ;
 wire \tms1x00.RAM[24][2] ;
 wire \tms1x00.RAM[24][3] ;
 wire \tms1x00.RAM[25][0] ;
 wire \tms1x00.RAM[25][1] ;
 wire \tms1x00.RAM[25][2] ;
 wire \tms1x00.RAM[25][3] ;
 wire \tms1x00.RAM[26][0] ;
 wire \tms1x00.RAM[26][1] ;
 wire \tms1x00.RAM[26][2] ;
 wire \tms1x00.RAM[26][3] ;
 wire \tms1x00.RAM[27][0] ;
 wire \tms1x00.RAM[27][1] ;
 wire \tms1x00.RAM[27][2] ;
 wire \tms1x00.RAM[27][3] ;
 wire \tms1x00.RAM[28][0] ;
 wire \tms1x00.RAM[28][1] ;
 wire \tms1x00.RAM[28][2] ;
 wire \tms1x00.RAM[28][3] ;
 wire \tms1x00.RAM[29][0] ;
 wire \tms1x00.RAM[29][1] ;
 wire \tms1x00.RAM[29][2] ;
 wire \tms1x00.RAM[29][3] ;
 wire \tms1x00.RAM[2][0] ;
 wire \tms1x00.RAM[2][1] ;
 wire \tms1x00.RAM[2][2] ;
 wire \tms1x00.RAM[2][3] ;
 wire \tms1x00.RAM[30][0] ;
 wire \tms1x00.RAM[30][1] ;
 wire \tms1x00.RAM[30][2] ;
 wire \tms1x00.RAM[30][3] ;
 wire \tms1x00.RAM[31][0] ;
 wire \tms1x00.RAM[31][1] ;
 wire \tms1x00.RAM[31][2] ;
 wire \tms1x00.RAM[31][3] ;
 wire \tms1x00.RAM[32][0] ;
 wire \tms1x00.RAM[32][1] ;
 wire \tms1x00.RAM[32][2] ;
 wire \tms1x00.RAM[32][3] ;
 wire \tms1x00.RAM[33][0] ;
 wire \tms1x00.RAM[33][1] ;
 wire \tms1x00.RAM[33][2] ;
 wire \tms1x00.RAM[33][3] ;
 wire \tms1x00.RAM[34][0] ;
 wire \tms1x00.RAM[34][1] ;
 wire \tms1x00.RAM[34][2] ;
 wire \tms1x00.RAM[34][3] ;
 wire \tms1x00.RAM[35][0] ;
 wire \tms1x00.RAM[35][1] ;
 wire \tms1x00.RAM[35][2] ;
 wire \tms1x00.RAM[35][3] ;
 wire \tms1x00.RAM[36][0] ;
 wire \tms1x00.RAM[36][1] ;
 wire \tms1x00.RAM[36][2] ;
 wire \tms1x00.RAM[36][3] ;
 wire \tms1x00.RAM[37][0] ;
 wire \tms1x00.RAM[37][1] ;
 wire \tms1x00.RAM[37][2] ;
 wire \tms1x00.RAM[37][3] ;
 wire \tms1x00.RAM[38][0] ;
 wire \tms1x00.RAM[38][1] ;
 wire \tms1x00.RAM[38][2] ;
 wire \tms1x00.RAM[38][3] ;
 wire \tms1x00.RAM[39][0] ;
 wire \tms1x00.RAM[39][1] ;
 wire \tms1x00.RAM[39][2] ;
 wire \tms1x00.RAM[39][3] ;
 wire \tms1x00.RAM[3][0] ;
 wire \tms1x00.RAM[3][1] ;
 wire \tms1x00.RAM[3][2] ;
 wire \tms1x00.RAM[3][3] ;
 wire \tms1x00.RAM[40][0] ;
 wire \tms1x00.RAM[40][1] ;
 wire \tms1x00.RAM[40][2] ;
 wire \tms1x00.RAM[40][3] ;
 wire \tms1x00.RAM[41][0] ;
 wire \tms1x00.RAM[41][1] ;
 wire \tms1x00.RAM[41][2] ;
 wire \tms1x00.RAM[41][3] ;
 wire \tms1x00.RAM[42][0] ;
 wire \tms1x00.RAM[42][1] ;
 wire \tms1x00.RAM[42][2] ;
 wire \tms1x00.RAM[42][3] ;
 wire \tms1x00.RAM[43][0] ;
 wire \tms1x00.RAM[43][1] ;
 wire \tms1x00.RAM[43][2] ;
 wire \tms1x00.RAM[43][3] ;
 wire \tms1x00.RAM[44][0] ;
 wire \tms1x00.RAM[44][1] ;
 wire \tms1x00.RAM[44][2] ;
 wire \tms1x00.RAM[44][3] ;
 wire \tms1x00.RAM[45][0] ;
 wire \tms1x00.RAM[45][1] ;
 wire \tms1x00.RAM[45][2] ;
 wire \tms1x00.RAM[45][3] ;
 wire \tms1x00.RAM[46][0] ;
 wire \tms1x00.RAM[46][1] ;
 wire \tms1x00.RAM[46][2] ;
 wire \tms1x00.RAM[46][3] ;
 wire \tms1x00.RAM[47][0] ;
 wire \tms1x00.RAM[47][1] ;
 wire \tms1x00.RAM[47][2] ;
 wire \tms1x00.RAM[47][3] ;
 wire \tms1x00.RAM[48][0] ;
 wire \tms1x00.RAM[48][1] ;
 wire \tms1x00.RAM[48][2] ;
 wire \tms1x00.RAM[48][3] ;
 wire \tms1x00.RAM[49][0] ;
 wire \tms1x00.RAM[49][1] ;
 wire \tms1x00.RAM[49][2] ;
 wire \tms1x00.RAM[49][3] ;
 wire \tms1x00.RAM[4][0] ;
 wire \tms1x00.RAM[4][1] ;
 wire \tms1x00.RAM[4][2] ;
 wire \tms1x00.RAM[4][3] ;
 wire \tms1x00.RAM[50][0] ;
 wire \tms1x00.RAM[50][1] ;
 wire \tms1x00.RAM[50][2] ;
 wire \tms1x00.RAM[50][3] ;
 wire \tms1x00.RAM[51][0] ;
 wire \tms1x00.RAM[51][1] ;
 wire \tms1x00.RAM[51][2] ;
 wire \tms1x00.RAM[51][3] ;
 wire \tms1x00.RAM[52][0] ;
 wire \tms1x00.RAM[52][1] ;
 wire \tms1x00.RAM[52][2] ;
 wire \tms1x00.RAM[52][3] ;
 wire \tms1x00.RAM[53][0] ;
 wire \tms1x00.RAM[53][1] ;
 wire \tms1x00.RAM[53][2] ;
 wire \tms1x00.RAM[53][3] ;
 wire \tms1x00.RAM[54][0] ;
 wire \tms1x00.RAM[54][1] ;
 wire \tms1x00.RAM[54][2] ;
 wire \tms1x00.RAM[54][3] ;
 wire \tms1x00.RAM[55][0] ;
 wire \tms1x00.RAM[55][1] ;
 wire \tms1x00.RAM[55][2] ;
 wire \tms1x00.RAM[55][3] ;
 wire \tms1x00.RAM[56][0] ;
 wire \tms1x00.RAM[56][1] ;
 wire \tms1x00.RAM[56][2] ;
 wire \tms1x00.RAM[56][3] ;
 wire \tms1x00.RAM[57][0] ;
 wire \tms1x00.RAM[57][1] ;
 wire \tms1x00.RAM[57][2] ;
 wire \tms1x00.RAM[57][3] ;
 wire \tms1x00.RAM[58][0] ;
 wire \tms1x00.RAM[58][1] ;
 wire \tms1x00.RAM[58][2] ;
 wire \tms1x00.RAM[58][3] ;
 wire \tms1x00.RAM[59][0] ;
 wire \tms1x00.RAM[59][1] ;
 wire \tms1x00.RAM[59][2] ;
 wire \tms1x00.RAM[59][3] ;
 wire \tms1x00.RAM[5][0] ;
 wire \tms1x00.RAM[5][1] ;
 wire \tms1x00.RAM[5][2] ;
 wire \tms1x00.RAM[5][3] ;
 wire \tms1x00.RAM[60][0] ;
 wire \tms1x00.RAM[60][1] ;
 wire \tms1x00.RAM[60][2] ;
 wire \tms1x00.RAM[60][3] ;
 wire \tms1x00.RAM[61][0] ;
 wire \tms1x00.RAM[61][1] ;
 wire \tms1x00.RAM[61][2] ;
 wire \tms1x00.RAM[61][3] ;
 wire \tms1x00.RAM[62][0] ;
 wire \tms1x00.RAM[62][1] ;
 wire \tms1x00.RAM[62][2] ;
 wire \tms1x00.RAM[62][3] ;
 wire \tms1x00.RAM[63][0] ;
 wire \tms1x00.RAM[63][1] ;
 wire \tms1x00.RAM[63][2] ;
 wire \tms1x00.RAM[63][3] ;
 wire \tms1x00.RAM[64][0] ;
 wire \tms1x00.RAM[64][1] ;
 wire \tms1x00.RAM[64][2] ;
 wire \tms1x00.RAM[64][3] ;
 wire \tms1x00.RAM[65][0] ;
 wire \tms1x00.RAM[65][1] ;
 wire \tms1x00.RAM[65][2] ;
 wire \tms1x00.RAM[65][3] ;
 wire \tms1x00.RAM[66][0] ;
 wire \tms1x00.RAM[66][1] ;
 wire \tms1x00.RAM[66][2] ;
 wire \tms1x00.RAM[66][3] ;
 wire \tms1x00.RAM[67][0] ;
 wire \tms1x00.RAM[67][1] ;
 wire \tms1x00.RAM[67][2] ;
 wire \tms1x00.RAM[67][3] ;
 wire \tms1x00.RAM[68][0] ;
 wire \tms1x00.RAM[68][1] ;
 wire \tms1x00.RAM[68][2] ;
 wire \tms1x00.RAM[68][3] ;
 wire \tms1x00.RAM[69][0] ;
 wire \tms1x00.RAM[69][1] ;
 wire \tms1x00.RAM[69][2] ;
 wire \tms1x00.RAM[69][3] ;
 wire \tms1x00.RAM[6][0] ;
 wire \tms1x00.RAM[6][1] ;
 wire \tms1x00.RAM[6][2] ;
 wire \tms1x00.RAM[6][3] ;
 wire \tms1x00.RAM[70][0] ;
 wire \tms1x00.RAM[70][1] ;
 wire \tms1x00.RAM[70][2] ;
 wire \tms1x00.RAM[70][3] ;
 wire \tms1x00.RAM[71][0] ;
 wire \tms1x00.RAM[71][1] ;
 wire \tms1x00.RAM[71][2] ;
 wire \tms1x00.RAM[71][3] ;
 wire \tms1x00.RAM[72][0] ;
 wire \tms1x00.RAM[72][1] ;
 wire \tms1x00.RAM[72][2] ;
 wire \tms1x00.RAM[72][3] ;
 wire \tms1x00.RAM[73][0] ;
 wire \tms1x00.RAM[73][1] ;
 wire \tms1x00.RAM[73][2] ;
 wire \tms1x00.RAM[73][3] ;
 wire \tms1x00.RAM[74][0] ;
 wire \tms1x00.RAM[74][1] ;
 wire \tms1x00.RAM[74][2] ;
 wire \tms1x00.RAM[74][3] ;
 wire \tms1x00.RAM[75][0] ;
 wire \tms1x00.RAM[75][1] ;
 wire \tms1x00.RAM[75][2] ;
 wire \tms1x00.RAM[75][3] ;
 wire \tms1x00.RAM[76][0] ;
 wire \tms1x00.RAM[76][1] ;
 wire \tms1x00.RAM[76][2] ;
 wire \tms1x00.RAM[76][3] ;
 wire \tms1x00.RAM[77][0] ;
 wire \tms1x00.RAM[77][1] ;
 wire \tms1x00.RAM[77][2] ;
 wire \tms1x00.RAM[77][3] ;
 wire \tms1x00.RAM[78][0] ;
 wire \tms1x00.RAM[78][1] ;
 wire \tms1x00.RAM[78][2] ;
 wire \tms1x00.RAM[78][3] ;
 wire \tms1x00.RAM[79][0] ;
 wire \tms1x00.RAM[79][1] ;
 wire \tms1x00.RAM[79][2] ;
 wire \tms1x00.RAM[79][3] ;
 wire \tms1x00.RAM[7][0] ;
 wire \tms1x00.RAM[7][1] ;
 wire \tms1x00.RAM[7][2] ;
 wire \tms1x00.RAM[7][3] ;
 wire \tms1x00.RAM[80][0] ;
 wire \tms1x00.RAM[80][1] ;
 wire \tms1x00.RAM[80][2] ;
 wire \tms1x00.RAM[80][3] ;
 wire \tms1x00.RAM[81][0] ;
 wire \tms1x00.RAM[81][1] ;
 wire \tms1x00.RAM[81][2] ;
 wire \tms1x00.RAM[81][3] ;
 wire \tms1x00.RAM[82][0] ;
 wire \tms1x00.RAM[82][1] ;
 wire \tms1x00.RAM[82][2] ;
 wire \tms1x00.RAM[82][3] ;
 wire \tms1x00.RAM[83][0] ;
 wire \tms1x00.RAM[83][1] ;
 wire \tms1x00.RAM[83][2] ;
 wire \tms1x00.RAM[83][3] ;
 wire \tms1x00.RAM[84][0] ;
 wire \tms1x00.RAM[84][1] ;
 wire \tms1x00.RAM[84][2] ;
 wire \tms1x00.RAM[84][3] ;
 wire \tms1x00.RAM[85][0] ;
 wire \tms1x00.RAM[85][1] ;
 wire \tms1x00.RAM[85][2] ;
 wire \tms1x00.RAM[85][3] ;
 wire \tms1x00.RAM[86][0] ;
 wire \tms1x00.RAM[86][1] ;
 wire \tms1x00.RAM[86][2] ;
 wire \tms1x00.RAM[86][3] ;
 wire \tms1x00.RAM[87][0] ;
 wire \tms1x00.RAM[87][1] ;
 wire \tms1x00.RAM[87][2] ;
 wire \tms1x00.RAM[87][3] ;
 wire \tms1x00.RAM[88][0] ;
 wire \tms1x00.RAM[88][1] ;
 wire \tms1x00.RAM[88][2] ;
 wire \tms1x00.RAM[88][3] ;
 wire \tms1x00.RAM[89][0] ;
 wire \tms1x00.RAM[89][1] ;
 wire \tms1x00.RAM[89][2] ;
 wire \tms1x00.RAM[89][3] ;
 wire \tms1x00.RAM[8][0] ;
 wire \tms1x00.RAM[8][1] ;
 wire \tms1x00.RAM[8][2] ;
 wire \tms1x00.RAM[8][3] ;
 wire \tms1x00.RAM[90][0] ;
 wire \tms1x00.RAM[90][1] ;
 wire \tms1x00.RAM[90][2] ;
 wire \tms1x00.RAM[90][3] ;
 wire \tms1x00.RAM[91][0] ;
 wire \tms1x00.RAM[91][1] ;
 wire \tms1x00.RAM[91][2] ;
 wire \tms1x00.RAM[91][3] ;
 wire \tms1x00.RAM[92][0] ;
 wire \tms1x00.RAM[92][1] ;
 wire \tms1x00.RAM[92][2] ;
 wire \tms1x00.RAM[92][3] ;
 wire \tms1x00.RAM[93][0] ;
 wire \tms1x00.RAM[93][1] ;
 wire \tms1x00.RAM[93][2] ;
 wire \tms1x00.RAM[93][3] ;
 wire \tms1x00.RAM[94][0] ;
 wire \tms1x00.RAM[94][1] ;
 wire \tms1x00.RAM[94][2] ;
 wire \tms1x00.RAM[94][3] ;
 wire \tms1x00.RAM[95][0] ;
 wire \tms1x00.RAM[95][1] ;
 wire \tms1x00.RAM[95][2] ;
 wire \tms1x00.RAM[95][3] ;
 wire \tms1x00.RAM[96][0] ;
 wire \tms1x00.RAM[96][1] ;
 wire \tms1x00.RAM[96][2] ;
 wire \tms1x00.RAM[96][3] ;
 wire \tms1x00.RAM[97][0] ;
 wire \tms1x00.RAM[97][1] ;
 wire \tms1x00.RAM[97][2] ;
 wire \tms1x00.RAM[97][3] ;
 wire \tms1x00.RAM[98][0] ;
 wire \tms1x00.RAM[98][1] ;
 wire \tms1x00.RAM[98][2] ;
 wire \tms1x00.RAM[98][3] ;
 wire \tms1x00.RAM[99][0] ;
 wire \tms1x00.RAM[99][1] ;
 wire \tms1x00.RAM[99][2] ;
 wire \tms1x00.RAM[99][3] ;
 wire \tms1x00.RAM[9][0] ;
 wire \tms1x00.RAM[9][1] ;
 wire \tms1x00.RAM[9][2] ;
 wire \tms1x00.RAM[9][3] ;
 wire \tms1x00.SR[0] ;
 wire \tms1x00.SR[1] ;
 wire \tms1x00.SR[2] ;
 wire \tms1x00.SR[3] ;
 wire \tms1x00.SR[4] ;
 wire \tms1x00.SR[5] ;
 wire \tms1x00.X[0] ;
 wire \tms1x00.X[1] ;
 wire \tms1x00.X[2] ;
 wire \tms1x00.Y[0] ;
 wire \tms1x00.Y[1] ;
 wire \tms1x00.Y[2] ;
 wire \tms1x00.Y[3] ;
 wire \tms1x00.ins_in[0] ;
 wire \tms1x00.ins_in[1] ;
 wire \tms1x00.ins_in[2] ;
 wire \tms1x00.ins_in[3] ;
 wire \tms1x00.ins_in[4] ;
 wire \tms1x00.ins_in[5] ;
 wire \tms1x00.ins_in[6] ;
 wire \tms1x00.ins_in[7] ;
 wire \tms1x00.ram_addr_buff[0] ;
 wire \tms1x00.ram_addr_buff[1] ;
 wire \tms1x00.ram_addr_buff[2] ;
 wire \tms1x00.ram_addr_buff[3] ;
 wire \tms1x00.ram_addr_buff[4] ;
 wire \tms1x00.ram_addr_buff[5] ;
 wire \tms1x00.ram_addr_buff[6] ;
 wire \tms1x00.rom_addr[0] ;
 wire \tms1x00.rom_addr[1] ;
 wire \tms1x00.status ;
 wire \tms1x00.wb_step ;
 wire \tms1x00.wb_step_state ;
 wire valid;
 wire wb_rst_override;
 wire \wbs_o_buff[0] ;
 wire \wbs_o_buff[10] ;
 wire \wbs_o_buff[11] ;
 wire \wbs_o_buff[12] ;
 wire \wbs_o_buff[13] ;
 wire \wbs_o_buff[14] ;
 wire \wbs_o_buff[15] ;
 wire \wbs_o_buff[16] ;
 wire \wbs_o_buff[17] ;
 wire \wbs_o_buff[18] ;
 wire \wbs_o_buff[19] ;
 wire \wbs_o_buff[1] ;
 wire \wbs_o_buff[20] ;
 wire \wbs_o_buff[21] ;
 wire \wbs_o_buff[22] ;
 wire \wbs_o_buff[23] ;
 wire \wbs_o_buff[24] ;
 wire \wbs_o_buff[25] ;
 wire \wbs_o_buff[26] ;
 wire \wbs_o_buff[27] ;
 wire \wbs_o_buff[28] ;
 wire \wbs_o_buff[29] ;
 wire \wbs_o_buff[2] ;
 wire \wbs_o_buff[30] ;
 wire \wbs_o_buff[31] ;
 wire \wbs_o_buff[3] ;
 wire \wbs_o_buff[4] ;
 wire \wbs_o_buff[5] ;
 wire \wbs_o_buff[6] ;
 wire \wbs_o_buff[7] ;
 wire \wbs_o_buff[8] ;
 wire \wbs_o_buff[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0_0_wb_clk_i;
 wire clknet_1_1_0_wb_clk_i;
 wire clknet_2_0_0_wb_clk_i;
 wire clknet_2_1_0_wb_clk_i;
 wire clknet_2_2_0_wb_clk_i;
 wire clknet_2_3_0_wb_clk_i;
 wire net204;

 sky130_fd_sc_hd__and2_1 _2206_ (.A(net70),
    .B(net61),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_2 _2207_ (.A(_0658_),
    .X(valid));
 sky130_fd_sc_hd__clkbuf_4 _2208_ (.A(net52),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_1 _2209_ (.A0(net17),
    .A1(\wbs_o_buff[0] ),
    .S(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__clkbuf_1 _2210_ (.A(_0660_),
    .X(net119));
 sky130_fd_sc_hd__mux2_1 _2211_ (.A0(net28),
    .A1(\wbs_o_buff[1] ),
    .S(_0659_),
    .X(_0661_));
 sky130_fd_sc_hd__clkbuf_1 _2212_ (.A(_0661_),
    .X(net130));
 sky130_fd_sc_hd__mux2_1 _2213_ (.A0(net39),
    .A1(\wbs_o_buff[2] ),
    .S(_0659_),
    .X(_0662_));
 sky130_fd_sc_hd__clkbuf_1 _2214_ (.A(_0662_),
    .X(net141));
 sky130_fd_sc_hd__mux2_1 _2215_ (.A0(net42),
    .A1(\wbs_o_buff[3] ),
    .S(_0659_),
    .X(_0663_));
 sky130_fd_sc_hd__clkbuf_1 _2216_ (.A(_0663_),
    .X(net144));
 sky130_fd_sc_hd__mux2_1 _2217_ (.A0(net43),
    .A1(\wbs_o_buff[4] ),
    .S(_0659_),
    .X(_0664_));
 sky130_fd_sc_hd__clkbuf_1 _2218_ (.A(_0664_),
    .X(net145));
 sky130_fd_sc_hd__mux2_1 _2219_ (.A0(net44),
    .A1(\wbs_o_buff[5] ),
    .S(_0659_),
    .X(_0665_));
 sky130_fd_sc_hd__clkbuf_1 _2220_ (.A(_0665_),
    .X(net146));
 sky130_fd_sc_hd__mux2_1 _2221_ (.A0(net45),
    .A1(\wbs_o_buff[6] ),
    .S(_0659_),
    .X(_0666_));
 sky130_fd_sc_hd__clkbuf_1 _2222_ (.A(_0666_),
    .X(net147));
 sky130_fd_sc_hd__mux2_1 _2223_ (.A0(net46),
    .A1(\wbs_o_buff[7] ),
    .S(_0659_),
    .X(_0667_));
 sky130_fd_sc_hd__clkbuf_1 _2224_ (.A(_0667_),
    .X(net148));
 sky130_fd_sc_hd__mux2_1 _2225_ (.A0(net47),
    .A1(\wbs_o_buff[8] ),
    .S(_0659_),
    .X(_0668_));
 sky130_fd_sc_hd__clkbuf_1 _2226_ (.A(_0668_),
    .X(net149));
 sky130_fd_sc_hd__mux2_1 _2227_ (.A0(net48),
    .A1(\wbs_o_buff[9] ),
    .S(_0659_),
    .X(_0669_));
 sky130_fd_sc_hd__clkbuf_1 _2228_ (.A(_0669_),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 _2229_ (.A(net52),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _2230_ (.A0(net18),
    .A1(\wbs_o_buff[10] ),
    .S(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__clkbuf_1 _2231_ (.A(_0671_),
    .X(net120));
 sky130_fd_sc_hd__mux2_1 _2232_ (.A0(net19),
    .A1(\wbs_o_buff[11] ),
    .S(_0670_),
    .X(_0672_));
 sky130_fd_sc_hd__clkbuf_1 _2233_ (.A(_0672_),
    .X(net121));
 sky130_fd_sc_hd__mux2_1 _2234_ (.A0(net20),
    .A1(\wbs_o_buff[12] ),
    .S(_0670_),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_1 _2235_ (.A(_0673_),
    .X(net122));
 sky130_fd_sc_hd__mux2_1 _2236_ (.A0(net21),
    .A1(\wbs_o_buff[13] ),
    .S(_0670_),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_1 _2237_ (.A(_0674_),
    .X(net123));
 sky130_fd_sc_hd__mux2_1 _2238_ (.A0(net22),
    .A1(\wbs_o_buff[14] ),
    .S(_0670_),
    .X(_0675_));
 sky130_fd_sc_hd__clkbuf_1 _2239_ (.A(_0675_),
    .X(net124));
 sky130_fd_sc_hd__mux2_1 _2240_ (.A0(net23),
    .A1(\wbs_o_buff[15] ),
    .S(_0670_),
    .X(_0676_));
 sky130_fd_sc_hd__clkbuf_1 _2241_ (.A(_0676_),
    .X(net125));
 sky130_fd_sc_hd__mux2_1 _2242_ (.A0(net24),
    .A1(\wbs_o_buff[16] ),
    .S(_0670_),
    .X(_0677_));
 sky130_fd_sc_hd__clkbuf_1 _2243_ (.A(_0677_),
    .X(net126));
 sky130_fd_sc_hd__mux2_1 _2244_ (.A0(net25),
    .A1(\wbs_o_buff[17] ),
    .S(_0670_),
    .X(_0678_));
 sky130_fd_sc_hd__clkbuf_1 _2245_ (.A(_0678_),
    .X(net127));
 sky130_fd_sc_hd__mux2_1 _2246_ (.A0(net26),
    .A1(\wbs_o_buff[18] ),
    .S(_0670_),
    .X(_0679_));
 sky130_fd_sc_hd__clkbuf_1 _2247_ (.A(_0679_),
    .X(net128));
 sky130_fd_sc_hd__mux2_1 _2248_ (.A0(net27),
    .A1(\wbs_o_buff[19] ),
    .S(_0670_),
    .X(_0680_));
 sky130_fd_sc_hd__clkbuf_1 _2249_ (.A(_0680_),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 _2250_ (.A(net52),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _2251_ (.A0(net29),
    .A1(\wbs_o_buff[20] ),
    .S(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__clkbuf_1 _2252_ (.A(_0682_),
    .X(net131));
 sky130_fd_sc_hd__mux2_1 _2253_ (.A0(net30),
    .A1(\wbs_o_buff[21] ),
    .S(_0681_),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_1 _2254_ (.A(_0683_),
    .X(net132));
 sky130_fd_sc_hd__mux2_1 _2255_ (.A0(net31),
    .A1(\wbs_o_buff[22] ),
    .S(_0681_),
    .X(_0684_));
 sky130_fd_sc_hd__clkbuf_1 _2256_ (.A(_0684_),
    .X(net133));
 sky130_fd_sc_hd__mux2_1 _2257_ (.A0(net32),
    .A1(\wbs_o_buff[23] ),
    .S(_0681_),
    .X(_0685_));
 sky130_fd_sc_hd__clkbuf_1 _2258_ (.A(_0685_),
    .X(net134));
 sky130_fd_sc_hd__mux2_1 _2259_ (.A0(net33),
    .A1(\wbs_o_buff[24] ),
    .S(_0681_),
    .X(_0686_));
 sky130_fd_sc_hd__clkbuf_1 _2260_ (.A(_0686_),
    .X(net135));
 sky130_fd_sc_hd__mux2_1 _2261_ (.A0(net34),
    .A1(\wbs_o_buff[25] ),
    .S(_0681_),
    .X(_0687_));
 sky130_fd_sc_hd__clkbuf_1 _2262_ (.A(_0687_),
    .X(net136));
 sky130_fd_sc_hd__mux2_1 _2263_ (.A0(net35),
    .A1(\wbs_o_buff[26] ),
    .S(_0681_),
    .X(_0688_));
 sky130_fd_sc_hd__clkbuf_1 _2264_ (.A(_0688_),
    .X(net137));
 sky130_fd_sc_hd__mux2_1 _2265_ (.A0(net36),
    .A1(\wbs_o_buff[27] ),
    .S(_0681_),
    .X(_0689_));
 sky130_fd_sc_hd__clkbuf_1 _2266_ (.A(_0689_),
    .X(net138));
 sky130_fd_sc_hd__mux2_1 _2267_ (.A0(net37),
    .A1(\wbs_o_buff[28] ),
    .S(_0681_),
    .X(_0690_));
 sky130_fd_sc_hd__clkbuf_1 _2268_ (.A(_0690_),
    .X(net139));
 sky130_fd_sc_hd__mux2_1 _2269_ (.A0(net38),
    .A1(\wbs_o_buff[29] ),
    .S(_0681_),
    .X(_0691_));
 sky130_fd_sc_hd__clkbuf_1 _2270_ (.A(_0691_),
    .X(net140));
 sky130_fd_sc_hd__mux2_1 _2271_ (.A0(net40),
    .A1(\wbs_o_buff[30] ),
    .S(net52),
    .X(_0692_));
 sky130_fd_sc_hd__clkbuf_1 _2272_ (.A(_0692_),
    .X(net142));
 sky130_fd_sc_hd__mux2_1 _2273_ (.A0(net41),
    .A1(\wbs_o_buff[31] ),
    .S(net52),
    .X(_0693_));
 sky130_fd_sc_hd__clkbuf_1 _2274_ (.A(_0693_),
    .X(net143));
 sky130_fd_sc_hd__mux2_1 _2275_ (.A0(net2),
    .A1(\K_override[0] ),
    .S(net152),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_1 _2276_ (.A(_0694_),
    .X(\tms1x00.K_in[0] ));
 sky130_fd_sc_hd__mux2_1 _2277_ (.A0(net3),
    .A1(\K_override[1] ),
    .S(net152),
    .X(_0695_));
 sky130_fd_sc_hd__clkbuf_1 _2278_ (.A(_0695_),
    .X(\tms1x00.K_in[1] ));
 sky130_fd_sc_hd__mux2_1 _2279_ (.A0(net4),
    .A1(\K_override[2] ),
    .S(net152),
    .X(_0696_));
 sky130_fd_sc_hd__clkbuf_1 _2280_ (.A(_0696_),
    .X(\tms1x00.K_in[2] ));
 sky130_fd_sc_hd__mux2_1 _2281_ (.A0(net5),
    .A1(\K_override[3] ),
    .S(net152),
    .X(_0697_));
 sky130_fd_sc_hd__clkbuf_1 _2282_ (.A(_0697_),
    .X(\tms1x00.K_in[3] ));
 sky130_fd_sc_hd__inv_2 _2283_ (.A(net71),
    .Y(net117));
 sky130_fd_sc_hd__and3_1 _2284_ (.A(net52),
    .B(net117),
    .C(valid),
    .X(_0698_));
 sky130_fd_sc_hd__buf_2 _2285_ (.A(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__buf_2 _2286_ (.A(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__nor2_2 _2287_ (.A(net49),
    .B(_0699_),
    .Y(_0701_));
 sky130_fd_sc_hd__buf_2 _2288_ (.A(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__a22o_1 _2289_ (.A1(net72),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\wbs_o_buff[0] ),
    .X(_0003_));
 sky130_fd_sc_hd__a22o_1 _2290_ (.A1(net73),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\wbs_o_buff[1] ),
    .X(_0014_));
 sky130_fd_sc_hd__a22o_1 _2291_ (.A1(net74),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\wbs_o_buff[2] ),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_1 _2292_ (.A1(net75),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\wbs_o_buff[3] ),
    .X(_0028_));
 sky130_fd_sc_hd__a22o_1 _2293_ (.A1(net76),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\wbs_o_buff[4] ),
    .X(_0029_));
 sky130_fd_sc_hd__a22o_1 _2294_ (.A1(net151),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\wbs_o_buff[5] ),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _2295_ (.A1(net78),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\wbs_o_buff[6] ),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_1 _2296_ (.A1(net79),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\wbs_o_buff[7] ),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_1 _2297_ (.A1(net80),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\wbs_o_buff[8] ),
    .X(_0033_));
 sky130_fd_sc_hd__a22o_1 _2298_ (.A1(net81),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\wbs_o_buff[9] ),
    .X(_0034_));
 sky130_fd_sc_hd__buf_2 _2299_ (.A(_0699_),
    .X(_0703_));
 sky130_fd_sc_hd__buf_2 _2300_ (.A(_0701_),
    .X(_0704_));
 sky130_fd_sc_hd__a22o_1 _2301_ (.A1(net82),
    .A2(_0703_),
    .B1(_0704_),
    .B2(\wbs_o_buff[10] ),
    .X(_0004_));
 sky130_fd_sc_hd__a22o_1 _2302_ (.A1(net83),
    .A2(_0703_),
    .B1(_0704_),
    .B2(\wbs_o_buff[11] ),
    .X(_0005_));
 sky130_fd_sc_hd__a22o_1 _2303_ (.A1(net84),
    .A2(_0703_),
    .B1(_0704_),
    .B2(\wbs_o_buff[12] ),
    .X(_0006_));
 sky130_fd_sc_hd__a22o_1 _2304_ (.A1(net85),
    .A2(_0703_),
    .B1(_0704_),
    .B2(\wbs_o_buff[13] ),
    .X(_0007_));
 sky130_fd_sc_hd__a22o_1 _2305_ (.A1(net86),
    .A2(_0703_),
    .B1(_0704_),
    .B2(\wbs_o_buff[14] ),
    .X(_0008_));
 sky130_fd_sc_hd__a22o_1 _2306_ (.A1(net87),
    .A2(_0703_),
    .B1(_0704_),
    .B2(\wbs_o_buff[15] ),
    .X(_0009_));
 sky130_fd_sc_hd__a22o_1 _2307_ (.A1(net88),
    .A2(_0703_),
    .B1(_0704_),
    .B2(\wbs_o_buff[16] ),
    .X(_0010_));
 sky130_fd_sc_hd__a22o_1 _2308_ (.A1(net89),
    .A2(_0703_),
    .B1(_0704_),
    .B2(\wbs_o_buff[17] ),
    .X(_0011_));
 sky130_fd_sc_hd__a22o_1 _2309_ (.A1(net90),
    .A2(_0703_),
    .B1(_0704_),
    .B2(\wbs_o_buff[18] ),
    .X(_0012_));
 sky130_fd_sc_hd__a22o_1 _2310_ (.A1(net91),
    .A2(_0703_),
    .B1(_0704_),
    .B2(\wbs_o_buff[19] ),
    .X(_0013_));
 sky130_fd_sc_hd__buf_2 _2311_ (.A(_0701_),
    .X(_0705_));
 sky130_fd_sc_hd__a22o_1 _2312_ (.A1(net92),
    .A2(_0699_),
    .B1(_0705_),
    .B2(\wbs_o_buff[20] ),
    .X(_0015_));
 sky130_fd_sc_hd__a22o_1 _2313_ (.A1(net93),
    .A2(_0699_),
    .B1(_0705_),
    .B2(\wbs_o_buff[21] ),
    .X(_0016_));
 sky130_fd_sc_hd__a22o_1 _2314_ (.A1(net94),
    .A2(_0699_),
    .B1(_0705_),
    .B2(\wbs_o_buff[22] ),
    .X(_0017_));
 sky130_fd_sc_hd__a22o_1 _2315_ (.A1(net95),
    .A2(_0699_),
    .B1(_0705_),
    .B2(\wbs_o_buff[23] ),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _2316_ (.A(\wbs_o_buff[24] ),
    .B(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__clkbuf_1 _2317_ (.A(_0706_),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _2318_ (.A(\wbs_o_buff[25] ),
    .B(_0705_),
    .X(_0707_));
 sky130_fd_sc_hd__clkbuf_1 _2319_ (.A(_0707_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _2320_ (.A(\wbs_o_buff[26] ),
    .B(_0705_),
    .X(_0708_));
 sky130_fd_sc_hd__clkbuf_1 _2321_ (.A(_0708_),
    .X(_0021_));
 sky130_fd_sc_hd__and2_1 _2322_ (.A(\wbs_o_buff[27] ),
    .B(_0705_),
    .X(_0709_));
 sky130_fd_sc_hd__clkbuf_1 _2323_ (.A(_0709_),
    .X(_0022_));
 sky130_fd_sc_hd__and2_1 _2324_ (.A(\wbs_o_buff[28] ),
    .B(_0705_),
    .X(_0710_));
 sky130_fd_sc_hd__clkbuf_1 _2325_ (.A(_0710_),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _2326_ (.A(\wbs_o_buff[29] ),
    .B(_0705_),
    .X(_0711_));
 sky130_fd_sc_hd__clkbuf_1 _2327_ (.A(_0711_),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _2328_ (.A(\wbs_o_buff[30] ),
    .B(_0701_),
    .X(_0712_));
 sky130_fd_sc_hd__clkbuf_1 _2329_ (.A(_0712_),
    .X(_0026_));
 sky130_fd_sc_hd__and2_1 _2330_ (.A(\wbs_o_buff[31] ),
    .B(_0701_),
    .X(_0713_));
 sky130_fd_sc_hd__clkbuf_1 _2331_ (.A(_0713_),
    .X(_0027_));
 sky130_fd_sc_hd__inv_2 _2332_ (.A(net49),
    .Y(_0714_));
 sky130_fd_sc_hd__nand3_2 _2333_ (.A(net52),
    .B(net71),
    .C(valid),
    .Y(_0715_));
 sky130_fd_sc_hd__and3_2 _2334_ (.A(net52),
    .B(net71),
    .C(valid),
    .X(_0716_));
 sky130_fd_sc_hd__and2_1 _2335_ (.A(net62),
    .B(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__a32o_1 _2336_ (.A1(wb_rst_override),
    .A2(_0714_),
    .A3(_0715_),
    .B1(_0717_),
    .B2(net65),
    .X(_0001_));
 sky130_fd_sc_hd__a32o_1 _2337_ (.A1(\tms1x00.wb_step ),
    .A2(_0714_),
    .A3(_0715_),
    .B1(_0717_),
    .B2(net66),
    .X(_0002_));
 sky130_fd_sc_hd__a31o_1 _2338_ (.A1(_0714_),
    .A2(net152),
    .A3(_0715_),
    .B1(_0717_),
    .X(_0000_));
 sky130_fd_sc_hd__nor2_4 _2339_ (.A(wb_rst_override),
    .B(net49),
    .Y(_0718_));
 sky130_fd_sc_hd__inv_2 _2340_ (.A(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__clkbuf_4 _2341_ (.A(_0719_),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 _2342_ (.A(\tms1x00.ram_addr_buff[0] ),
    .X(_0720_));
 sky130_fd_sc_hd__or3b_2 _2343_ (.A(net78),
    .B(net151),
    .C_N(net79),
    .X(_0721_));
 sky130_fd_sc_hd__xnor2_2 _2344_ (.A(\tms1x00.wb_step ),
    .B(\tms1x00.wb_step_state ),
    .Y(_0722_));
 sky130_fd_sc_hd__a21o_1 _2345_ (.A1(net152),
    .A2(_0722_),
    .B1(_0719_),
    .X(_0723_));
 sky130_fd_sc_hd__or2_2 _2346_ (.A(_0721_),
    .B(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__clkbuf_4 _2347_ (.A(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _2348_ (.A0(\tms1x00.Y[0] ),
    .A1(_0720_),
    .S(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__clkbuf_1 _2349_ (.A(_0726_),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_2 _2350_ (.A(\tms1x00.ram_addr_buff[1] ),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _2351_ (.A0(\tms1x00.Y[1] ),
    .A1(_0727_),
    .S(_0725_),
    .X(_0728_));
 sky130_fd_sc_hd__clkbuf_1 _2352_ (.A(_0728_),
    .X(_0043_));
 sky130_fd_sc_hd__buf_2 _2353_ (.A(\tms1x00.Y[2] ),
    .X(_0729_));
 sky130_fd_sc_hd__buf_2 _2354_ (.A(\tms1x00.ram_addr_buff[2] ),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _2355_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0725_),
    .X(_0731_));
 sky130_fd_sc_hd__clkbuf_1 _2356_ (.A(_0731_),
    .X(_0044_));
 sky130_fd_sc_hd__buf_2 _2357_ (.A(\tms1x00.Y[3] ),
    .X(_0732_));
 sky130_fd_sc_hd__buf_2 _2358_ (.A(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__buf_2 _2359_ (.A(\tms1x00.ram_addr_buff[3] ),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _2360_ (.A0(_0733_),
    .A1(_0734_),
    .S(_0725_),
    .X(_0735_));
 sky130_fd_sc_hd__clkbuf_1 _2361_ (.A(_0735_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2362_ (.A0(\tms1x00.X[2] ),
    .A1(\tms1x00.ram_addr_buff[4] ),
    .S(_0725_),
    .X(_0736_));
 sky130_fd_sc_hd__clkbuf_1 _2363_ (.A(_0736_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2364_ (.A0(\tms1x00.X[0] ),
    .A1(\tms1x00.ram_addr_buff[5] ),
    .S(_0725_),
    .X(_0737_));
 sky130_fd_sc_hd__clkbuf_1 _2365_ (.A(_0737_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _2366_ (.A0(\tms1x00.X[1] ),
    .A1(\tms1x00.ram_addr_buff[6] ),
    .S(_0725_),
    .X(_0738_));
 sky130_fd_sc_hd__clkbuf_1 _2367_ (.A(_0738_),
    .X(_0048_));
 sky130_fd_sc_hd__nand2_1 _2368_ (.A(net51),
    .B(valid),
    .Y(net116));
 sky130_fd_sc_hd__clkinv_2 _2369_ (.A(\tms1x00.Y[2] ),
    .Y(_0739_));
 sky130_fd_sc_hd__nor2_1 _2370_ (.A(\tms1x00.Y[1] ),
    .B(\tms1x00.Y[0] ),
    .Y(_0740_));
 sky130_fd_sc_hd__nand2_1 _2371_ (.A(_0739_),
    .B(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__clkbuf_4 _2372_ (.A(\tms1x00.ins_in[7] ),
    .X(_0742_));
 sky130_fd_sc_hd__buf_2 _2373_ (.A(\tms1x00.ins_in[4] ),
    .X(_0743_));
 sky130_fd_sc_hd__nand2_1 _2374_ (.A(\tms1x00.ins_in[5] ),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__and2_2 _2375_ (.A(net152),
    .B(_0722_),
    .X(_0745_));
 sky130_fd_sc_hd__nand3b_2 _2376_ (.A_N(net79),
    .B(net78),
    .C(net151),
    .Y(_0746_));
 sky130_fd_sc_hd__or2_1 _2377_ (.A(_0745_),
    .B(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__or4_1 _2378_ (.A(\tms1x00.ins_in[3] ),
    .B(\tms1x00.ins_in[2] ),
    .C(\tms1x00.ins_in[1] ),
    .D(\tms1x00.ins_in[0] ),
    .X(_0748_));
 sky130_fd_sc_hd__or2_1 _2379_ (.A(_0747_),
    .B(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__or4_4 _2380_ (.A(_0742_),
    .B(\tms1x00.ins_in[6] ),
    .C(_0744_),
    .D(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__buf_2 _2381_ (.A(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__inv_2 _2382_ (.A(\tms1x00.Y[3] ),
    .Y(_0752_));
 sky130_fd_sc_hd__buf_2 _2383_ (.A(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__and2_1 _2384_ (.A(_0739_),
    .B(_0740_),
    .X(_0754_));
 sky130_fd_sc_hd__clkinv_2 _2385_ (.A(_0742_),
    .Y(_0755_));
 sky130_fd_sc_hd__nor2_1 _2386_ (.A(_0755_),
    .B(\tms1x00.ins_in[6] ),
    .Y(_0756_));
 sky130_fd_sc_hd__a21oi_2 _2387_ (.A1(net152),
    .A2(_0722_),
    .B1(_0746_),
    .Y(_0757_));
 sky130_fd_sc_hd__nor2_1 _2388_ (.A(_0748_),
    .B(_0744_),
    .Y(_0758_));
 sky130_fd_sc_hd__and3_2 _2389_ (.A(_0756_),
    .B(_0757_),
    .C(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__buf_2 _2390_ (.A(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__a31o_1 _2391_ (.A1(_0753_),
    .A2(_0754_),
    .A3(_0760_),
    .B1(net80),
    .X(_0761_));
 sky130_fd_sc_hd__clkbuf_4 _2392_ (.A(_0718_),
    .X(_0762_));
 sky130_fd_sc_hd__o311a_1 _2393_ (.A1(_0733_),
    .A2(_0741_),
    .A3(_0751_),
    .B1(_0761_),
    .C1(_0762_),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_1 _2394_ (.A1(chip_sel_override),
    .A2(_0715_),
    .B1(_0717_),
    .B2(net67),
    .X(_0050_));
 sky130_fd_sc_hd__clkinv_2 _2395_ (.A(\tms1x00.ins_in[6] ),
    .Y(_0763_));
 sky130_fd_sc_hd__clkinv_2 _2396_ (.A(_0040_),
    .Y(_0764_));
 sky130_fd_sc_hd__clkinv_2 _2397_ (.A(_0038_),
    .Y(_0765_));
 sky130_fd_sc_hd__clkbuf_4 _2398_ (.A(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__clkbuf_4 _2399_ (.A(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__buf_8 _2400_ (.A(_0035_),
    .X(_0768_));
 sky130_fd_sc_hd__buf_8 _2401_ (.A(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__buf_6 _2402_ (.A(_0036_),
    .X(_0770_));
 sky130_fd_sc_hd__buf_8 _2403_ (.A(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__mux4_1 _2404_ (.A0(\tms1x00.RAM[80][0] ),
    .A1(\tms1x00.RAM[81][0] ),
    .A2(\tms1x00.RAM[82][0] ),
    .A3(\tms1x00.RAM[83][0] ),
    .S0(_0769_),
    .S1(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__buf_6 _2405_ (.A(_0035_),
    .X(_0773_));
 sky130_fd_sc_hd__buf_8 _2406_ (.A(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__mux4_1 _2407_ (.A0(\tms1x00.RAM[84][0] ),
    .A1(\tms1x00.RAM[85][0] ),
    .A2(\tms1x00.RAM[86][0] ),
    .A3(\tms1x00.RAM[87][0] ),
    .S0(_0774_),
    .S1(_0771_),
    .X(_0775_));
 sky130_fd_sc_hd__clkbuf_4 _2408_ (.A(_0037_),
    .X(_0776_));
 sky130_fd_sc_hd__buf_4 _2409_ (.A(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _2410_ (.A0(_0772_),
    .A1(_0775_),
    .S(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__buf_4 _2411_ (.A(_0036_),
    .X(_0779_));
 sky130_fd_sc_hd__buf_4 _2412_ (.A(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__buf_4 _2413_ (.A(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__buf_6 _2414_ (.A(_0035_),
    .X(_0782_));
 sky130_fd_sc_hd__mux2_1 _2415_ (.A0(\tms1x00.RAM[94][0] ),
    .A1(\tms1x00.RAM[95][0] ),
    .S(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__and2_1 _2416_ (.A(_0781_),
    .B(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__inv_2 _2417_ (.A(_0779_),
    .Y(_0785_));
 sky130_fd_sc_hd__buf_4 _2418_ (.A(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__buf_6 _2419_ (.A(_0035_),
    .X(_0787_));
 sky130_fd_sc_hd__mux2_1 _2420_ (.A0(\tms1x00.RAM[92][0] ),
    .A1(\tms1x00.RAM[93][0] ),
    .S(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__inv_2 _2421_ (.A(_0037_),
    .Y(_0789_));
 sky130_fd_sc_hd__buf_4 _2422_ (.A(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__a21o_1 _2423_ (.A1(_0786_),
    .A2(_0788_),
    .B1(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__buf_6 _2424_ (.A(_0770_),
    .X(_0792_));
 sky130_fd_sc_hd__mux4_1 _2425_ (.A0(\tms1x00.RAM[88][0] ),
    .A1(\tms1x00.RAM[89][0] ),
    .A2(\tms1x00.RAM[90][0] ),
    .A3(\tms1x00.RAM[91][0] ),
    .S0(_0769_),
    .S1(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__buf_4 _2426_ (.A(_0776_),
    .X(_0794_));
 sky130_fd_sc_hd__buf_4 _2427_ (.A(_0038_),
    .X(_0795_));
 sky130_fd_sc_hd__o221a_1 _2428_ (.A1(_0784_),
    .A2(_0791_),
    .B1(_0793_),
    .B2(_0794_),
    .C1(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__inv_2 _2429_ (.A(_0039_),
    .Y(_0797_));
 sky130_fd_sc_hd__clkbuf_4 _2430_ (.A(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__a211o_1 _2431_ (.A1(_0767_),
    .A2(_0778_),
    .B1(_0796_),
    .C1(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__clkbuf_4 _2432_ (.A(_0038_),
    .X(_0800_));
 sky130_fd_sc_hd__clkbuf_4 _2433_ (.A(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__clkbuf_4 _2434_ (.A(_0776_),
    .X(_0802_));
 sky130_fd_sc_hd__clkbuf_8 _2435_ (.A(_0773_),
    .X(_0803_));
 sky130_fd_sc_hd__buf_6 _2436_ (.A(_0779_),
    .X(_0804_));
 sky130_fd_sc_hd__mux4_1 _2437_ (.A0(\tms1x00.RAM[72][0] ),
    .A1(\tms1x00.RAM[73][0] ),
    .A2(\tms1x00.RAM[74][0] ),
    .A3(\tms1x00.RAM[75][0] ),
    .S0(_0803_),
    .S1(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__or2_1 _2438_ (.A(_0802_),
    .B(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__buf_4 _2439_ (.A(_0787_),
    .X(_0807_));
 sky130_fd_sc_hd__or2b_1 _2440_ (.A(\tms1x00.RAM[79][0] ),
    .B_N(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__clkbuf_4 _2441_ (.A(_0770_),
    .X(_0809_));
 sky130_fd_sc_hd__o21a_1 _2442_ (.A1(_0807_),
    .A2(\tms1x00.RAM[78][0] ),
    .B1(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__buf_6 _2443_ (.A(_0035_),
    .X(_0811_));
 sky130_fd_sc_hd__buf_6 _2444_ (.A(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _2445_ (.A0(\tms1x00.RAM[76][0] ),
    .A1(\tms1x00.RAM[77][0] ),
    .S(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__buf_4 _2446_ (.A(_0785_),
    .X(_0814_));
 sky130_fd_sc_hd__clkbuf_4 _2447_ (.A(_0789_),
    .X(_0815_));
 sky130_fd_sc_hd__buf_4 _2448_ (.A(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__a221o_1 _2449_ (.A1(_0808_),
    .A2(_0810_),
    .B1(_0813_),
    .B2(_0814_),
    .C1(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__clkbuf_4 _2450_ (.A(_0039_),
    .X(_0818_));
 sky130_fd_sc_hd__mux2_1 _2451_ (.A0(\tms1x00.RAM[70][0] ),
    .A1(\tms1x00.RAM[71][0] ),
    .S(_0782_),
    .X(_0819_));
 sky130_fd_sc_hd__and2_1 _2452_ (.A(_0809_),
    .B(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _2453_ (.A0(\tms1x00.RAM[68][0] ),
    .A1(\tms1x00.RAM[69][0] ),
    .S(_0787_),
    .X(_0821_));
 sky130_fd_sc_hd__a21o_1 _2454_ (.A1(_0786_),
    .A2(_0821_),
    .B1(_0815_),
    .X(_0822_));
 sky130_fd_sc_hd__mux4_2 _2455_ (.A0(\tms1x00.RAM[64][0] ),
    .A1(\tms1x00.RAM[65][0] ),
    .A2(\tms1x00.RAM[66][0] ),
    .A3(\tms1x00.RAM[67][0] ),
    .S0(_0774_),
    .S1(_0771_),
    .X(_0823_));
 sky130_fd_sc_hd__clkbuf_4 _2456_ (.A(_0765_),
    .X(_0824_));
 sky130_fd_sc_hd__o221a_1 _2457_ (.A1(_0820_),
    .A2(_0822_),
    .B1(_0823_),
    .B2(_0794_),
    .C1(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__a311o_1 _2458_ (.A1(_0801_),
    .A2(_0806_),
    .A3(_0817_),
    .B1(_0818_),
    .C1(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__inv_2 _2459_ (.A(_0041_),
    .Y(_0827_));
 sky130_fd_sc_hd__buf_4 _2460_ (.A(_0790_),
    .X(_0828_));
 sky130_fd_sc_hd__mux4_1 _2461_ (.A0(\tms1x00.RAM[108][0] ),
    .A1(\tms1x00.RAM[109][0] ),
    .A2(\tms1x00.RAM[110][0] ),
    .A3(\tms1x00.RAM[111][0] ),
    .S0(_0769_),
    .S1(_0792_),
    .X(_0829_));
 sky130_fd_sc_hd__mux4_1 _2462_ (.A0(\tms1x00.RAM[104][0] ),
    .A1(\tms1x00.RAM[105][0] ),
    .A2(\tms1x00.RAM[106][0] ),
    .A3(\tms1x00.RAM[107][0] ),
    .S0(_0773_),
    .S1(_0779_),
    .X(_0830_));
 sky130_fd_sc_hd__or2_1 _2463_ (.A(_0776_),
    .B(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__o211a_1 _2464_ (.A1(_0828_),
    .A2(_0829_),
    .B1(_0831_),
    .C1(_0795_),
    .X(_0832_));
 sky130_fd_sc_hd__buf_6 _2465_ (.A(_0768_),
    .X(_0833_));
 sky130_fd_sc_hd__mux4_1 _2466_ (.A0(\tms1x00.RAM[96][0] ),
    .A1(\tms1x00.RAM[97][0] ),
    .A2(\tms1x00.RAM[98][0] ),
    .A3(\tms1x00.RAM[99][0] ),
    .S0(_0833_),
    .S1(_0809_),
    .X(_0834_));
 sky130_fd_sc_hd__mux4_1 _2467_ (.A0(\tms1x00.RAM[100][0] ),
    .A1(\tms1x00.RAM[101][0] ),
    .A2(\tms1x00.RAM[102][0] ),
    .A3(\tms1x00.RAM[103][0] ),
    .S0(_0768_),
    .S1(_0770_),
    .X(_0835_));
 sky130_fd_sc_hd__or2_1 _2468_ (.A(_0790_),
    .B(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__o211a_1 _2469_ (.A1(_0794_),
    .A2(_0834_),
    .B1(_0836_),
    .C1(_0824_),
    .X(_0837_));
 sky130_fd_sc_hd__mux4_1 _2470_ (.A0(\tms1x00.RAM[120][0] ),
    .A1(\tms1x00.RAM[121][0] ),
    .A2(\tms1x00.RAM[122][0] ),
    .A3(\tms1x00.RAM[123][0] ),
    .S0(_0768_),
    .S1(_0770_),
    .X(_0838_));
 sky130_fd_sc_hd__or2_1 _2471_ (.A(_0776_),
    .B(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__buf_4 _2472_ (.A(_0036_),
    .X(_0840_));
 sky130_fd_sc_hd__mux4_1 _2473_ (.A0(\tms1x00.RAM[124][0] ),
    .A1(\tms1x00.RAM[125][0] ),
    .A2(\tms1x00.RAM[126][0] ),
    .A3(\tms1x00.RAM[127][0] ),
    .S0(_0811_),
    .S1(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__o21a_1 _2474_ (.A1(_0790_),
    .A2(_0841_),
    .B1(_0038_),
    .X(_0842_));
 sky130_fd_sc_hd__or2b_1 _2475_ (.A(\tms1x00.RAM[119][0] ),
    .B_N(_0803_),
    .X(_0843_));
 sky130_fd_sc_hd__buf_6 _2476_ (.A(_0773_),
    .X(_0844_));
 sky130_fd_sc_hd__o21a_1 _2477_ (.A1(_0844_),
    .A2(\tms1x00.RAM[118][0] ),
    .B1(_0780_),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_1 _2478_ (.A0(\tms1x00.RAM[116][0] ),
    .A1(\tms1x00.RAM[117][0] ),
    .S(_0787_),
    .X(_0846_));
 sky130_fd_sc_hd__a221o_1 _2479_ (.A1(_0843_),
    .A2(_0845_),
    .B1(_0846_),
    .B2(_0786_),
    .C1(_0790_),
    .X(_0847_));
 sky130_fd_sc_hd__buf_4 _2480_ (.A(_0776_),
    .X(_0848_));
 sky130_fd_sc_hd__mux4_1 _2481_ (.A0(\tms1x00.RAM[112][0] ),
    .A1(\tms1x00.RAM[113][0] ),
    .A2(\tms1x00.RAM[114][0] ),
    .A3(\tms1x00.RAM[115][0] ),
    .S0(_0811_),
    .S1(_0840_),
    .X(_0849_));
 sky130_fd_sc_hd__o21a_1 _2482_ (.A1(_0848_),
    .A2(_0849_),
    .B1(_0765_),
    .X(_0850_));
 sky130_fd_sc_hd__a221o_1 _2483_ (.A1(_0839_),
    .A2(_0842_),
    .B1(_0847_),
    .B2(_0850_),
    .C1(_0797_),
    .X(_0851_));
 sky130_fd_sc_hd__o311a_1 _2484_ (.A1(_0818_),
    .A2(_0832_),
    .A3(_0837_),
    .B1(_0851_),
    .C1(_0040_),
    .X(_0852_));
 sky130_fd_sc_hd__a311o_2 _2485_ (.A1(_0764_),
    .A2(_0799_),
    .A3(_0826_),
    .B1(_0827_),
    .C1(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__mux4_1 _2486_ (.A0(\tms1x00.RAM[16][0] ),
    .A1(\tms1x00.RAM[17][0] ),
    .A2(\tms1x00.RAM[18][0] ),
    .A3(\tms1x00.RAM[19][0] ),
    .S0(_0769_),
    .S1(_0792_),
    .X(_0854_));
 sky130_fd_sc_hd__mux4_1 _2487_ (.A0(\tms1x00.RAM[20][0] ),
    .A1(\tms1x00.RAM[21][0] ),
    .A2(\tms1x00.RAM[22][0] ),
    .A3(\tms1x00.RAM[23][0] ),
    .S0(_0769_),
    .S1(_0771_),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _2488_ (.A0(_0854_),
    .A1(_0855_),
    .S(_0802_),
    .X(_0856_));
 sky130_fd_sc_hd__clkbuf_4 _2489_ (.A(_0785_),
    .X(_0857_));
 sky130_fd_sc_hd__buf_6 _2490_ (.A(_0844_),
    .X(_0858_));
 sky130_fd_sc_hd__mux2_1 _2491_ (.A0(\tms1x00.RAM[28][0] ),
    .A1(\tms1x00.RAM[29][0] ),
    .S(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__buf_6 _2492_ (.A(_0804_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _2493_ (.A0(\tms1x00.RAM[30][0] ),
    .A1(\tms1x00.RAM[31][0] ),
    .S(_0774_),
    .X(_0861_));
 sky130_fd_sc_hd__buf_4 _2494_ (.A(_0815_),
    .X(_0862_));
 sky130_fd_sc_hd__a21o_1 _2495_ (.A1(_0860_),
    .A2(_0861_),
    .B1(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__a21o_1 _2496_ (.A1(_0857_),
    .A2(_0859_),
    .B1(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__buf_4 _2497_ (.A(_0848_),
    .X(_0865_));
 sky130_fd_sc_hd__mux4_1 _2498_ (.A0(\tms1x00.RAM[24][0] ),
    .A1(\tms1x00.RAM[25][0] ),
    .A2(\tms1x00.RAM[26][0] ),
    .A3(\tms1x00.RAM[27][0] ),
    .S0(_0812_),
    .S1(_0781_),
    .X(_0866_));
 sky130_fd_sc_hd__o21a_1 _2499_ (.A1(_0865_),
    .A2(_0866_),
    .B1(_0795_),
    .X(_0867_));
 sky130_fd_sc_hd__a221o_1 _2500_ (.A1(_0767_),
    .A2(_0856_),
    .B1(_0864_),
    .B2(_0867_),
    .C1(_0798_),
    .X(_0868_));
 sky130_fd_sc_hd__mux4_1 _2501_ (.A0(\tms1x00.RAM[8][0] ),
    .A1(\tms1x00.RAM[9][0] ),
    .A2(\tms1x00.RAM[10][0] ),
    .A3(\tms1x00.RAM[11][0] ),
    .S0(_0833_),
    .S1(_0792_),
    .X(_0869_));
 sky130_fd_sc_hd__or2_1 _2502_ (.A(_0794_),
    .B(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__or2b_1 _2503_ (.A(\tms1x00.RAM[15][0] ),
    .B_N(_0858_),
    .X(_0871_));
 sky130_fd_sc_hd__o21a_1 _2504_ (.A1(_0858_),
    .A2(\tms1x00.RAM[14][0] ),
    .B1(_0781_),
    .X(_0872_));
 sky130_fd_sc_hd__buf_4 _2505_ (.A(_0782_),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(\tms1x00.RAM[12][0] ),
    .A1(\tms1x00.RAM[13][0] ),
    .S(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__a221o_1 _2507_ (.A1(_0871_),
    .A2(_0872_),
    .B1(_0874_),
    .B2(_0857_),
    .C1(_0828_),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _2508_ (.A0(\tms1x00.RAM[6][0] ),
    .A1(\tms1x00.RAM[7][0] ),
    .S(_0787_),
    .X(_0876_));
 sky130_fd_sc_hd__and2_1 _2509_ (.A(_0781_),
    .B(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(\tms1x00.RAM[4][0] ),
    .A1(\tms1x00.RAM[5][0] ),
    .S(_0787_),
    .X(_0878_));
 sky130_fd_sc_hd__a21o_1 _2511_ (.A1(_0786_),
    .A2(_0878_),
    .B1(_0862_),
    .X(_0879_));
 sky130_fd_sc_hd__mux4_1 _2512_ (.A0(\tms1x00.RAM[0][0] ),
    .A1(\tms1x00.RAM[1][0] ),
    .A2(\tms1x00.RAM[2][0] ),
    .A3(\tms1x00.RAM[3][0] ),
    .S0(_0833_),
    .S1(_0809_),
    .X(_0880_));
 sky130_fd_sc_hd__o221a_1 _2513_ (.A1(_0877_),
    .A2(_0879_),
    .B1(_0880_),
    .B2(_0865_),
    .C1(_0824_),
    .X(_0881_));
 sky130_fd_sc_hd__a311o_1 _2514_ (.A1(_0801_),
    .A2(_0870_),
    .A3(_0875_),
    .B1(_0818_),
    .C1(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__mux4_1 _2515_ (.A0(\tms1x00.RAM[44][0] ),
    .A1(\tms1x00.RAM[45][0] ),
    .A2(\tms1x00.RAM[46][0] ),
    .A3(\tms1x00.RAM[47][0] ),
    .S0(_0768_),
    .S1(_0840_),
    .X(_0883_));
 sky130_fd_sc_hd__or2_1 _2516_ (.A(_0790_),
    .B(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__mux4_1 _2517_ (.A0(\tms1x00.RAM[40][0] ),
    .A1(\tms1x00.RAM[41][0] ),
    .A2(\tms1x00.RAM[42][0] ),
    .A3(\tms1x00.RAM[43][0] ),
    .S0(_0811_),
    .S1(_0840_),
    .X(_0885_));
 sky130_fd_sc_hd__o21a_1 _2518_ (.A1(_0848_),
    .A2(_0885_),
    .B1(_0800_),
    .X(_0886_));
 sky130_fd_sc_hd__mux4_1 _2519_ (.A0(\tms1x00.RAM[32][0] ),
    .A1(\tms1x00.RAM[33][0] ),
    .A2(\tms1x00.RAM[34][0] ),
    .A3(\tms1x00.RAM[35][0] ),
    .S0(_0811_),
    .S1(_0840_),
    .X(_0887_));
 sky130_fd_sc_hd__or2_1 _2520_ (.A(_0848_),
    .B(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__mux4_2 _2521_ (.A0(\tms1x00.RAM[36][0] ),
    .A1(\tms1x00.RAM[37][0] ),
    .A2(\tms1x00.RAM[38][0] ),
    .A3(\tms1x00.RAM[39][0] ),
    .S0(_0811_),
    .S1(_0840_),
    .X(_0889_));
 sky130_fd_sc_hd__o21a_1 _2522_ (.A1(_0862_),
    .A2(_0889_),
    .B1(_0766_),
    .X(_0890_));
 sky130_fd_sc_hd__a221o_1 _2523_ (.A1(_0884_),
    .A2(_0886_),
    .B1(_0888_),
    .B2(_0890_),
    .C1(_0039_),
    .X(_0891_));
 sky130_fd_sc_hd__mux4_1 _2524_ (.A0(\tms1x00.RAM[56][0] ),
    .A1(\tms1x00.RAM[57][0] ),
    .A2(\tms1x00.RAM[58][0] ),
    .A3(\tms1x00.RAM[59][0] ),
    .S0(_0768_),
    .S1(_0770_),
    .X(_0892_));
 sky130_fd_sc_hd__or2_1 _2525_ (.A(_0848_),
    .B(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__mux4_2 _2526_ (.A0(\tms1x00.RAM[60][0] ),
    .A1(\tms1x00.RAM[61][0] ),
    .A2(\tms1x00.RAM[62][0] ),
    .A3(\tms1x00.RAM[63][0] ),
    .S0(_0811_),
    .S1(_0840_),
    .X(_0894_));
 sky130_fd_sc_hd__o21a_1 _2527_ (.A1(_0862_),
    .A2(_0894_),
    .B1(_0800_),
    .X(_0895_));
 sky130_fd_sc_hd__or2b_1 _2528_ (.A(\tms1x00.RAM[55][0] ),
    .B_N(_0803_),
    .X(_0896_));
 sky130_fd_sc_hd__o21a_1 _2529_ (.A1(_0803_),
    .A2(\tms1x00.RAM[54][0] ),
    .B1(_0780_),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(\tms1x00.RAM[52][0] ),
    .A1(\tms1x00.RAM[53][0] ),
    .S(_0787_),
    .X(_0898_));
 sky130_fd_sc_hd__a221o_1 _2531_ (.A1(_0896_),
    .A2(_0897_),
    .B1(_0898_),
    .B2(_0786_),
    .C1(_0790_),
    .X(_0899_));
 sky130_fd_sc_hd__mux4_1 _2532_ (.A0(\tms1x00.RAM[48][0] ),
    .A1(\tms1x00.RAM[49][0] ),
    .A2(\tms1x00.RAM[50][0] ),
    .A3(\tms1x00.RAM[51][0] ),
    .S0(_0811_),
    .S1(_0840_),
    .X(_0900_));
 sky130_fd_sc_hd__o21a_1 _2533_ (.A1(_0848_),
    .A2(_0900_),
    .B1(_0766_),
    .X(_0901_));
 sky130_fd_sc_hd__a221o_1 _2534_ (.A1(_0893_),
    .A2(_0895_),
    .B1(_0899_),
    .B2(_0901_),
    .C1(_0797_),
    .X(_0902_));
 sky130_fd_sc_hd__a31o_1 _2535_ (.A1(_0040_),
    .A2(_0891_),
    .A3(_0902_),
    .B1(_0041_),
    .X(_0903_));
 sky130_fd_sc_hd__a31o_2 _2536_ (.A1(_0764_),
    .A2(_0868_),
    .A3(_0882_),
    .B1(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__a22o_1 _2537_ (.A1(_0755_),
    .A2(_0763_),
    .B1(_0853_),
    .B2(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__nor2_1 _2538_ (.A(\tms1x00.ins_in[1] ),
    .B(\tms1x00.ins_in[0] ),
    .Y(_0906_));
 sky130_fd_sc_hd__and3_1 _2539_ (.A(\tms1x00.ins_in[3] ),
    .B(\tms1x00.ins_in[2] ),
    .C(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__and4b_1 _2540_ (.A_N(\tms1x00.ins_in[4] ),
    .B(_0718_),
    .C(_0757_),
    .D(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__or2b_1 _2541_ (.A(\tms1x00.ins_in[5] ),
    .B_N(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__inv_2 _2542_ (.A(\tms1x00.ins_in[3] ),
    .Y(_0910_));
 sky130_fd_sc_hd__and4b_1 _2543_ (.A_N(\tms1x00.ins_in[5] ),
    .B(\tms1x00.ins_in[4] ),
    .C(\tms1x00.ins_in[7] ),
    .D(\tms1x00.ins_in[6] ),
    .X(_0911_));
 sky130_fd_sc_hd__nand3_1 _2544_ (.A(_0910_),
    .B(\tms1x00.ins_in[2] ),
    .C(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__or4b_1 _2545_ (.A(net79),
    .B(net151),
    .C(\tms1x00.ins_in[1] ),
    .D_N(net78),
    .X(_0913_));
 sky130_fd_sc_hd__nor3_2 _2546_ (.A(_0723_),
    .B(_0912_),
    .C(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__a31oi_1 _2547_ (.A1(_0755_),
    .A2(_0763_),
    .A3(_0909_),
    .B1(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__nor3_2 _2548_ (.A(_0723_),
    .B(_0912_),
    .C(_0913_),
    .Y(_0916_));
 sky130_fd_sc_hd__and3_1 _2549_ (.A(\tms1x00.A[0] ),
    .B(_0906_),
    .C(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__a21o_1 _2550_ (.A1(_0905_),
    .A2(_0915_),
    .B1(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__buf_4 _2551_ (.A(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__clkbuf_4 _2552_ (.A(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__nand3b_2 _2553_ (.A_N(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[6] ),
    .Y(_0921_));
 sky130_fd_sc_hd__buf_4 _2554_ (.A(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__or2b_2 _2555_ (.A(_0727_),
    .B_N(_0720_),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_1 _2556_ (.A(\tms1x00.ram_addr_buff[2] ),
    .B(\tms1x00.ram_addr_buff[3] ),
    .Y(_0924_));
 sky130_fd_sc_hd__nor2_1 _2557_ (.A(\tms1x00.ins_in[4] ),
    .B(_0747_),
    .Y(_0925_));
 sky130_fd_sc_hd__a31oi_4 _2558_ (.A1(_0718_),
    .A2(_0925_),
    .A3(_0907_),
    .B1(_0914_),
    .Y(_0926_));
 sky130_fd_sc_hd__or3_1 _2559_ (.A(_0923_),
    .B(_0924_),
    .C(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__buf_6 _2560_ (.A(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__nor2_2 _2561_ (.A(_0922_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__mux2_1 _2562_ (.A0(\tms1x00.RAM[109][0] ),
    .A1(_0920_),
    .S(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__clkbuf_1 _2563_ (.A(_0930_),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _2564_ (.A(_0906_),
    .B(_0916_),
    .X(_0931_));
 sky130_fd_sc_hd__buf_8 _2565_ (.A(_0773_),
    .X(_0932_));
 sky130_fd_sc_hd__buf_6 _2566_ (.A(_0779_),
    .X(_0933_));
 sky130_fd_sc_hd__mux4_1 _2567_ (.A0(\tms1x00.RAM[80][1] ),
    .A1(\tms1x00.RAM[81][1] ),
    .A2(\tms1x00.RAM[82][1] ),
    .A3(\tms1x00.RAM[83][1] ),
    .S0(_0932_),
    .S1(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__mux4_1 _2568_ (.A0(\tms1x00.RAM[84][1] ),
    .A1(\tms1x00.RAM[85][1] ),
    .A2(\tms1x00.RAM[86][1] ),
    .A3(\tms1x00.RAM[87][1] ),
    .S0(_0932_),
    .S1(_0933_),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(_0934_),
    .A1(_0935_),
    .S(_0848_),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_1 _2570_ (.A0(\tms1x00.RAM[92][1] ),
    .A1(\tms1x00.RAM[93][1] ),
    .S(_0807_),
    .X(_0937_));
 sky130_fd_sc_hd__clkbuf_8 _2571_ (.A(_0780_),
    .X(_0938_));
 sky130_fd_sc_hd__buf_6 _2572_ (.A(_0773_),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(\tms1x00.RAM[94][1] ),
    .A1(\tms1x00.RAM[95][1] ),
    .S(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__a21o_1 _2574_ (.A1(_0938_),
    .A2(_0940_),
    .B1(_0862_),
    .X(_0941_));
 sky130_fd_sc_hd__a21o_1 _2575_ (.A1(_0857_),
    .A2(_0937_),
    .B1(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__mux4_1 _2576_ (.A0(\tms1x00.RAM[88][1] ),
    .A1(\tms1x00.RAM[89][1] ),
    .A2(\tms1x00.RAM[90][1] ),
    .A3(\tms1x00.RAM[91][1] ),
    .S0(_0833_),
    .S1(_0792_),
    .X(_0943_));
 sky130_fd_sc_hd__o21a_1 _2577_ (.A1(_0794_),
    .A2(_0943_),
    .B1(_0795_),
    .X(_0944_));
 sky130_fd_sc_hd__a221o_1 _2578_ (.A1(_0767_),
    .A2(_0936_),
    .B1(_0942_),
    .B2(_0944_),
    .C1(_0798_),
    .X(_0945_));
 sky130_fd_sc_hd__buf_6 _2579_ (.A(_0779_),
    .X(_0946_));
 sky130_fd_sc_hd__mux4_1 _2580_ (.A0(\tms1x00.RAM[72][1] ),
    .A1(\tms1x00.RAM[73][1] ),
    .A2(\tms1x00.RAM[74][1] ),
    .A3(\tms1x00.RAM[75][1] ),
    .S0(_0844_),
    .S1(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__or2_1 _2581_ (.A(_0802_),
    .B(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__or2b_1 _2582_ (.A(\tms1x00.RAM[79][1] ),
    .B_N(_0807_),
    .X(_0949_));
 sky130_fd_sc_hd__o21a_1 _2583_ (.A1(_0807_),
    .A2(\tms1x00.RAM[78][1] ),
    .B1(_0809_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _2584_ (.A0(\tms1x00.RAM[76][1] ),
    .A1(\tms1x00.RAM[77][1] ),
    .S(_0812_),
    .X(_0951_));
 sky130_fd_sc_hd__a221o_1 _2585_ (.A1(_0949_),
    .A2(_0950_),
    .B1(_0951_),
    .B2(_0814_),
    .C1(_0816_),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_1 _2586_ (.A0(\tms1x00.RAM[70][1] ),
    .A1(\tms1x00.RAM[71][1] ),
    .S(_0782_),
    .X(_0953_));
 sky130_fd_sc_hd__and2_1 _2587_ (.A(_0809_),
    .B(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__mux2_1 _2588_ (.A0(\tms1x00.RAM[68][1] ),
    .A1(\tms1x00.RAM[69][1] ),
    .S(_0782_),
    .X(_0955_));
 sky130_fd_sc_hd__a21o_1 _2589_ (.A1(_0786_),
    .A2(_0955_),
    .B1(_0815_),
    .X(_0956_));
 sky130_fd_sc_hd__mux4_2 _2590_ (.A0(\tms1x00.RAM[64][1] ),
    .A1(\tms1x00.RAM[65][1] ),
    .A2(\tms1x00.RAM[66][1] ),
    .A3(\tms1x00.RAM[67][1] ),
    .S0(_0774_),
    .S1(_0771_),
    .X(_0957_));
 sky130_fd_sc_hd__o221a_1 _2591_ (.A1(_0954_),
    .A2(_0956_),
    .B1(_0957_),
    .B2(_0794_),
    .C1(_0824_),
    .X(_0958_));
 sky130_fd_sc_hd__a311o_1 _2592_ (.A1(_0801_),
    .A2(_0948_),
    .A3(_0952_),
    .B1(_0818_),
    .C1(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__mux4_1 _2593_ (.A0(\tms1x00.RAM[108][1] ),
    .A1(\tms1x00.RAM[109][1] ),
    .A2(\tms1x00.RAM[110][1] ),
    .A3(\tms1x00.RAM[111][1] ),
    .S0(_0769_),
    .S1(_0792_),
    .X(_0960_));
 sky130_fd_sc_hd__mux4_1 _2594_ (.A0(\tms1x00.RAM[104][1] ),
    .A1(\tms1x00.RAM[105][1] ),
    .A2(\tms1x00.RAM[106][1] ),
    .A3(\tms1x00.RAM[107][1] ),
    .S0(_0773_),
    .S1(_0779_),
    .X(_0961_));
 sky130_fd_sc_hd__or2_1 _2595_ (.A(_0776_),
    .B(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__o211a_1 _2596_ (.A1(_0828_),
    .A2(_0960_),
    .B1(_0962_),
    .C1(_0795_),
    .X(_0963_));
 sky130_fd_sc_hd__mux4_1 _2597_ (.A0(\tms1x00.RAM[96][1] ),
    .A1(\tms1x00.RAM[97][1] ),
    .A2(\tms1x00.RAM[98][1] ),
    .A3(\tms1x00.RAM[99][1] ),
    .S0(_0833_),
    .S1(_0809_),
    .X(_0964_));
 sky130_fd_sc_hd__mux4_1 _2598_ (.A0(\tms1x00.RAM[100][1] ),
    .A1(\tms1x00.RAM[101][1] ),
    .A2(\tms1x00.RAM[102][1] ),
    .A3(\tms1x00.RAM[103][1] ),
    .S0(_0768_),
    .S1(_0770_),
    .X(_0965_));
 sky130_fd_sc_hd__or2_1 _2599_ (.A(_0790_),
    .B(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__o211a_1 _2600_ (.A1(_0794_),
    .A2(_0964_),
    .B1(_0966_),
    .C1(_0824_),
    .X(_0967_));
 sky130_fd_sc_hd__mux4_1 _2601_ (.A0(\tms1x00.RAM[120][1] ),
    .A1(\tms1x00.RAM[121][1] ),
    .A2(\tms1x00.RAM[122][1] ),
    .A3(\tms1x00.RAM[123][1] ),
    .S0(_0768_),
    .S1(_0770_),
    .X(_0968_));
 sky130_fd_sc_hd__or2_1 _2602_ (.A(_0776_),
    .B(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__mux4_1 _2603_ (.A0(\tms1x00.RAM[124][1] ),
    .A1(\tms1x00.RAM[125][1] ),
    .A2(\tms1x00.RAM[126][1] ),
    .A3(\tms1x00.RAM[127][1] ),
    .S0(_0811_),
    .S1(_0840_),
    .X(_0970_));
 sky130_fd_sc_hd__o21a_1 _2604_ (.A1(_0790_),
    .A2(_0970_),
    .B1(_0038_),
    .X(_0971_));
 sky130_fd_sc_hd__or2b_1 _2605_ (.A(\tms1x00.RAM[119][1] ),
    .B_N(_0844_),
    .X(_0972_));
 sky130_fd_sc_hd__o21a_1 _2606_ (.A1(_0844_),
    .A2(\tms1x00.RAM[118][1] ),
    .B1(_0780_),
    .X(_0973_));
 sky130_fd_sc_hd__mux2_1 _2607_ (.A0(\tms1x00.RAM[116][1] ),
    .A1(\tms1x00.RAM[117][1] ),
    .S(_0787_),
    .X(_0974_));
 sky130_fd_sc_hd__a221o_1 _2608_ (.A1(_0972_),
    .A2(_0973_),
    .B1(_0974_),
    .B2(_0786_),
    .C1(_0790_),
    .X(_0975_));
 sky130_fd_sc_hd__mux4_1 _2609_ (.A0(\tms1x00.RAM[112][1] ),
    .A1(\tms1x00.RAM[113][1] ),
    .A2(\tms1x00.RAM[114][1] ),
    .A3(\tms1x00.RAM[115][1] ),
    .S0(_0811_),
    .S1(_0840_),
    .X(_0976_));
 sky130_fd_sc_hd__o21a_1 _2610_ (.A1(_0848_),
    .A2(_0976_),
    .B1(_0765_),
    .X(_0977_));
 sky130_fd_sc_hd__a221o_1 _2611_ (.A1(_0969_),
    .A2(_0971_),
    .B1(_0975_),
    .B2(_0977_),
    .C1(_0797_),
    .X(_0978_));
 sky130_fd_sc_hd__o311a_1 _2612_ (.A1(_0818_),
    .A2(_0963_),
    .A3(_0967_),
    .B1(_0978_),
    .C1(_0040_),
    .X(_0979_));
 sky130_fd_sc_hd__a311o_1 _2613_ (.A1(_0764_),
    .A2(_0945_),
    .A3(_0959_),
    .B1(_0827_),
    .C1(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__mux4_1 _2614_ (.A0(\tms1x00.RAM[16][1] ),
    .A1(\tms1x00.RAM[17][1] ),
    .A2(\tms1x00.RAM[18][1] ),
    .A3(\tms1x00.RAM[19][1] ),
    .S0(_0774_),
    .S1(_0771_),
    .X(_0981_));
 sky130_fd_sc_hd__mux4_2 _2615_ (.A0(\tms1x00.RAM[20][1] ),
    .A1(\tms1x00.RAM[21][1] ),
    .A2(\tms1x00.RAM[22][1] ),
    .A3(\tms1x00.RAM[23][1] ),
    .S0(_0774_),
    .S1(_0804_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _2616_ (.A0(_0981_),
    .A1(_0982_),
    .S(_0777_),
    .X(_0983_));
 sky130_fd_sc_hd__mux2_1 _2617_ (.A0(\tms1x00.RAM[30][1] ),
    .A1(\tms1x00.RAM[31][1] ),
    .S(_0782_),
    .X(_0984_));
 sky130_fd_sc_hd__and2_1 _2618_ (.A(_0809_),
    .B(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _2619_ (.A0(\tms1x00.RAM[28][1] ),
    .A1(\tms1x00.RAM[29][1] ),
    .S(_0782_),
    .X(_0986_));
 sky130_fd_sc_hd__a21o_1 _2620_ (.A1(_0786_),
    .A2(_0986_),
    .B1(_0815_),
    .X(_0987_));
 sky130_fd_sc_hd__mux4_2 _2621_ (.A0(\tms1x00.RAM[24][1] ),
    .A1(\tms1x00.RAM[25][1] ),
    .A2(\tms1x00.RAM[26][1] ),
    .A3(\tms1x00.RAM[27][1] ),
    .S0(_0774_),
    .S1(_0771_),
    .X(_0988_));
 sky130_fd_sc_hd__o221a_1 _2622_ (.A1(_0985_),
    .A2(_0987_),
    .B1(_0988_),
    .B2(_0794_),
    .C1(_0795_),
    .X(_0989_));
 sky130_fd_sc_hd__a211o_1 _2623_ (.A1(_0767_),
    .A2(_0983_),
    .B1(_0989_),
    .C1(_0798_),
    .X(_0990_));
 sky130_fd_sc_hd__mux4_1 _2624_ (.A0(\tms1x00.RAM[8][1] ),
    .A1(\tms1x00.RAM[9][1] ),
    .A2(\tms1x00.RAM[10][1] ),
    .A3(\tms1x00.RAM[11][1] ),
    .S0(_0932_),
    .S1(_0946_),
    .X(_0991_));
 sky130_fd_sc_hd__or2_1 _2625_ (.A(_0802_),
    .B(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__or2b_1 _2626_ (.A(\tms1x00.RAM[15][1] ),
    .B_N(_0807_),
    .X(_0993_));
 sky130_fd_sc_hd__buf_4 _2627_ (.A(_0787_),
    .X(_0994_));
 sky130_fd_sc_hd__o21a_1 _2628_ (.A1(_0994_),
    .A2(\tms1x00.RAM[14][1] ),
    .B1(_0792_),
    .X(_0995_));
 sky130_fd_sc_hd__mux2_1 _2629_ (.A0(\tms1x00.RAM[12][1] ),
    .A1(\tms1x00.RAM[13][1] ),
    .S(_0812_),
    .X(_0996_));
 sky130_fd_sc_hd__clkbuf_4 _2630_ (.A(_0815_),
    .X(_0997_));
 sky130_fd_sc_hd__a221o_1 _2631_ (.A1(_0993_),
    .A2(_0995_),
    .B1(_0996_),
    .B2(_0814_),
    .C1(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(\tms1x00.RAM[6][1] ),
    .A1(\tms1x00.RAM[7][1] ),
    .S(_0782_),
    .X(_0999_));
 sky130_fd_sc_hd__and2_1 _2633_ (.A(_0809_),
    .B(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(\tms1x00.RAM[4][1] ),
    .A1(\tms1x00.RAM[5][1] ),
    .S(_0782_),
    .X(_1001_));
 sky130_fd_sc_hd__a21o_1 _2635_ (.A1(_0785_),
    .A2(_1001_),
    .B1(_0815_),
    .X(_1002_));
 sky130_fd_sc_hd__mux4_1 _2636_ (.A0(\tms1x00.RAM[0][1] ),
    .A1(\tms1x00.RAM[1][1] ),
    .A2(\tms1x00.RAM[2][1] ),
    .A3(\tms1x00.RAM[3][1] ),
    .S0(_0803_),
    .S1(_0804_),
    .X(_1003_));
 sky130_fd_sc_hd__o221a_1 _2637_ (.A1(_1000_),
    .A2(_1002_),
    .B1(_1003_),
    .B2(_0802_),
    .C1(_0766_),
    .X(_1004_));
 sky130_fd_sc_hd__a311o_1 _2638_ (.A1(_0801_),
    .A2(_0992_),
    .A3(_0998_),
    .B1(_0039_),
    .C1(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__mux4_1 _2639_ (.A0(\tms1x00.RAM[44][1] ),
    .A1(\tms1x00.RAM[45][1] ),
    .A2(\tms1x00.RAM[46][1] ),
    .A3(\tms1x00.RAM[47][1] ),
    .S0(_0803_),
    .S1(_0804_),
    .X(_1006_));
 sky130_fd_sc_hd__mux4_1 _2640_ (.A0(\tms1x00.RAM[40][1] ),
    .A1(\tms1x00.RAM[41][1] ),
    .A2(\tms1x00.RAM[42][1] ),
    .A3(\tms1x00.RAM[43][1] ),
    .S0(_0773_),
    .S1(_0779_),
    .X(_1007_));
 sky130_fd_sc_hd__or2_1 _2641_ (.A(_0776_),
    .B(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__o211a_1 _2642_ (.A1(_0816_),
    .A2(_1006_),
    .B1(_1008_),
    .C1(_0800_),
    .X(_1009_));
 sky130_fd_sc_hd__mux4_1 _2643_ (.A0(\tms1x00.RAM[32][1] ),
    .A1(\tms1x00.RAM[33][1] ),
    .A2(\tms1x00.RAM[34][1] ),
    .A3(\tms1x00.RAM[35][1] ),
    .S0(_0769_),
    .S1(_0771_),
    .X(_1010_));
 sky130_fd_sc_hd__mux4_1 _2644_ (.A0(\tms1x00.RAM[36][1] ),
    .A1(\tms1x00.RAM[37][1] ),
    .A2(\tms1x00.RAM[38][1] ),
    .A3(\tms1x00.RAM[39][1] ),
    .S0(_0773_),
    .S1(_0779_),
    .X(_1011_));
 sky130_fd_sc_hd__or2_1 _2645_ (.A(_0815_),
    .B(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__o211a_1 _2646_ (.A1(_0794_),
    .A2(_1010_),
    .B1(_1012_),
    .C1(_0824_),
    .X(_1013_));
 sky130_fd_sc_hd__mux4_1 _2647_ (.A0(\tms1x00.RAM[56][1] ),
    .A1(\tms1x00.RAM[57][1] ),
    .A2(\tms1x00.RAM[58][1] ),
    .A3(\tms1x00.RAM[59][1] ),
    .S0(_0773_),
    .S1(_0779_),
    .X(_1014_));
 sky130_fd_sc_hd__or2_1 _2648_ (.A(_0776_),
    .B(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__mux4_2 _2649_ (.A0(\tms1x00.RAM[60][1] ),
    .A1(\tms1x00.RAM[61][1] ),
    .A2(\tms1x00.RAM[62][1] ),
    .A3(\tms1x00.RAM[63][1] ),
    .S0(_0768_),
    .S1(_0770_),
    .X(_1016_));
 sky130_fd_sc_hd__o21a_1 _2650_ (.A1(_0815_),
    .A2(_1016_),
    .B1(_0038_),
    .X(_1017_));
 sky130_fd_sc_hd__or2b_1 _2651_ (.A(\tms1x00.RAM[55][1] ),
    .B_N(_0939_),
    .X(_1018_));
 sky130_fd_sc_hd__o21a_1 _2652_ (.A1(_0939_),
    .A2(\tms1x00.RAM[54][1] ),
    .B1(_0780_),
    .X(_1019_));
 sky130_fd_sc_hd__mux2_1 _2653_ (.A0(\tms1x00.RAM[52][1] ),
    .A1(\tms1x00.RAM[53][1] ),
    .S(_0782_),
    .X(_1020_));
 sky130_fd_sc_hd__a221o_1 _2654_ (.A1(_1018_),
    .A2(_1019_),
    .B1(_1020_),
    .B2(_0785_),
    .C1(_0815_),
    .X(_1021_));
 sky130_fd_sc_hd__mux4_2 _2655_ (.A0(\tms1x00.RAM[48][1] ),
    .A1(\tms1x00.RAM[49][1] ),
    .A2(\tms1x00.RAM[50][1] ),
    .A3(\tms1x00.RAM[51][1] ),
    .S0(_0768_),
    .S1(_0770_),
    .X(_1022_));
 sky130_fd_sc_hd__o21a_1 _2656_ (.A1(_0848_),
    .A2(_1022_),
    .B1(_0765_),
    .X(_1023_));
 sky130_fd_sc_hd__a221o_1 _2657_ (.A1(_1015_),
    .A2(_1017_),
    .B1(_1021_),
    .B2(_1023_),
    .C1(_0797_),
    .X(_1024_));
 sky130_fd_sc_hd__o311a_1 _2658_ (.A1(_0039_),
    .A2(_1009_),
    .A3(_1013_),
    .B1(_1024_),
    .C1(_0040_),
    .X(_1025_));
 sky130_fd_sc_hd__a311o_2 _2659_ (.A1(_0764_),
    .A2(_0990_),
    .A3(_1005_),
    .B1(_1025_),
    .C1(_0041_),
    .X(_1026_));
 sky130_fd_sc_hd__nor2_2 _2660_ (.A(_0742_),
    .B(_0763_),
    .Y(_1027_));
 sky130_fd_sc_hd__a21o_1 _2661_ (.A1(_0980_),
    .A2(_1026_),
    .B1(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__a21oi_1 _2662_ (.A1(_0909_),
    .A2(_1027_),
    .B1(_0914_),
    .Y(_1029_));
 sky130_fd_sc_hd__a22o_2 _2663_ (.A1(\tms1x00.A[1] ),
    .A2(_0931_),
    .B1(_1028_),
    .B2(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__buf_4 _2664_ (.A(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__clkbuf_4 _2665_ (.A(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__mux2_1 _2666_ (.A0(\tms1x00.RAM[109][1] ),
    .A1(_1032_),
    .S(_0929_),
    .X(_1033_));
 sky130_fd_sc_hd__clkbuf_1 _2667_ (.A(_1033_),
    .X(_0052_));
 sky130_fd_sc_hd__mux4_1 _2668_ (.A0(\tms1x00.RAM[80][2] ),
    .A1(\tms1x00.RAM[81][2] ),
    .A2(\tms1x00.RAM[82][2] ),
    .A3(\tms1x00.RAM[83][2] ),
    .S0(_0858_),
    .S1(_0860_),
    .X(_1034_));
 sky130_fd_sc_hd__mux4_1 _2669_ (.A0(\tms1x00.RAM[84][2] ),
    .A1(\tms1x00.RAM[85][2] ),
    .A2(\tms1x00.RAM[86][2] ),
    .A3(\tms1x00.RAM[87][2] ),
    .S0(_0858_),
    .S1(_0860_),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _2670_ (.A0(_1034_),
    .A1(_1035_),
    .S(_0865_),
    .X(_1036_));
 sky130_fd_sc_hd__clkbuf_4 _2671_ (.A(_0780_),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _2672_ (.A0(\tms1x00.RAM[94][2] ),
    .A1(\tms1x00.RAM[95][2] ),
    .S(_0812_),
    .X(_1038_));
 sky130_fd_sc_hd__and2_1 _2673_ (.A(_1037_),
    .B(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _2674_ (.A0(\tms1x00.RAM[92][2] ),
    .A1(\tms1x00.RAM[93][2] ),
    .S(_0873_),
    .X(_1040_));
 sky130_fd_sc_hd__a21o_1 _2675_ (.A1(_0857_),
    .A2(_1040_),
    .B1(_0816_),
    .X(_1041_));
 sky130_fd_sc_hd__buf_4 _2676_ (.A(_0774_),
    .X(_1042_));
 sky130_fd_sc_hd__mux4_1 _2677_ (.A0(\tms1x00.RAM[88][2] ),
    .A1(\tms1x00.RAM[89][2] ),
    .A2(\tms1x00.RAM[90][2] ),
    .A3(\tms1x00.RAM[91][2] ),
    .S0(_1042_),
    .S1(_1037_),
    .X(_1043_));
 sky130_fd_sc_hd__clkbuf_4 _2678_ (.A(_0777_),
    .X(_1044_));
 sky130_fd_sc_hd__o221a_1 _2679_ (.A1(_1039_),
    .A2(_1041_),
    .B1(_1043_),
    .B2(_1044_),
    .C1(_0801_),
    .X(_1045_));
 sky130_fd_sc_hd__a211o_1 _2680_ (.A1(_0767_),
    .A2(_1036_),
    .B1(_1045_),
    .C1(_0798_),
    .X(_1046_));
 sky130_fd_sc_hd__buf_6 _2681_ (.A(_0939_),
    .X(_1047_));
 sky130_fd_sc_hd__mux4_1 _2682_ (.A0(\tms1x00.RAM[72][2] ),
    .A1(\tms1x00.RAM[73][2] ),
    .A2(\tms1x00.RAM[74][2] ),
    .A3(\tms1x00.RAM[75][2] ),
    .S0(_1047_),
    .S1(_0938_),
    .X(_1048_));
 sky130_fd_sc_hd__or2_1 _2683_ (.A(_1044_),
    .B(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__or2b_1 _2684_ (.A(\tms1x00.RAM[79][2] ),
    .B_N(_1042_),
    .X(_1050_));
 sky130_fd_sc_hd__o21a_1 _2685_ (.A1(_1042_),
    .A2(\tms1x00.RAM[78][2] ),
    .B1(_1037_),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_1 _2686_ (.A0(\tms1x00.RAM[76][2] ),
    .A1(\tms1x00.RAM[77][2] ),
    .S(_1042_),
    .X(_1052_));
 sky130_fd_sc_hd__a221o_1 _2687_ (.A1(_1050_),
    .A2(_1051_),
    .B1(_1052_),
    .B2(_0857_),
    .C1(_0828_),
    .X(_1053_));
 sky130_fd_sc_hd__mux2_1 _2688_ (.A0(\tms1x00.RAM[70][2] ),
    .A1(\tms1x00.RAM[71][2] ),
    .S(_0812_),
    .X(_1054_));
 sky130_fd_sc_hd__and2_1 _2689_ (.A(_1037_),
    .B(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__mux2_1 _2690_ (.A0(\tms1x00.RAM[68][2] ),
    .A1(\tms1x00.RAM[69][2] ),
    .S(_0812_),
    .X(_1056_));
 sky130_fd_sc_hd__a21o_1 _2691_ (.A1(_0857_),
    .A2(_1056_),
    .B1(_0816_),
    .X(_1057_));
 sky130_fd_sc_hd__mux4_1 _2692_ (.A0(\tms1x00.RAM[64][2] ),
    .A1(\tms1x00.RAM[65][2] ),
    .A2(\tms1x00.RAM[66][2] ),
    .A3(\tms1x00.RAM[67][2] ),
    .S0(_0858_),
    .S1(_0860_),
    .X(_1058_));
 sky130_fd_sc_hd__o221a_1 _2693_ (.A1(_1055_),
    .A2(_1057_),
    .B1(_1058_),
    .B2(_1044_),
    .C1(_0767_),
    .X(_1059_));
 sky130_fd_sc_hd__a311o_1 _2694_ (.A1(_0801_),
    .A2(_1049_),
    .A3(_1053_),
    .B1(_0818_),
    .C1(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__mux4_1 _2695_ (.A0(\tms1x00.RAM[120][2] ),
    .A1(\tms1x00.RAM[121][2] ),
    .A2(\tms1x00.RAM[122][2] ),
    .A3(\tms1x00.RAM[123][2] ),
    .S0(_0932_),
    .S1(_0933_),
    .X(_1061_));
 sky130_fd_sc_hd__or2_1 _2696_ (.A(_0777_),
    .B(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__mux4_1 _2697_ (.A0(\tms1x00.RAM[124][2] ),
    .A1(\tms1x00.RAM[125][2] ),
    .A2(\tms1x00.RAM[126][2] ),
    .A3(\tms1x00.RAM[127][2] ),
    .S0(_0844_),
    .S1(_0946_),
    .X(_1063_));
 sky130_fd_sc_hd__o21a_1 _2698_ (.A1(_0816_),
    .A2(_1063_),
    .B1(_0800_),
    .X(_1064_));
 sky130_fd_sc_hd__or2b_1 _2699_ (.A(\tms1x00.RAM[119][2] ),
    .B_N(_0994_),
    .X(_1065_));
 sky130_fd_sc_hd__o21a_1 _2700_ (.A1(_0994_),
    .A2(\tms1x00.RAM[118][2] ),
    .B1(_0792_),
    .X(_1066_));
 sky130_fd_sc_hd__mux2_1 _2701_ (.A0(\tms1x00.RAM[116][2] ),
    .A1(\tms1x00.RAM[117][2] ),
    .S(_0812_),
    .X(_1067_));
 sky130_fd_sc_hd__a221o_1 _2702_ (.A1(_1065_),
    .A2(_1066_),
    .B1(_1067_),
    .B2(_0814_),
    .C1(_0997_),
    .X(_1068_));
 sky130_fd_sc_hd__mux4_1 _2703_ (.A0(\tms1x00.RAM[112][2] ),
    .A1(\tms1x00.RAM[113][2] ),
    .A2(\tms1x00.RAM[114][2] ),
    .A3(\tms1x00.RAM[115][2] ),
    .S0(_0803_),
    .S1(_0804_),
    .X(_1069_));
 sky130_fd_sc_hd__o21a_1 _2704_ (.A1(_0802_),
    .A2(_1069_),
    .B1(_0766_),
    .X(_1070_));
 sky130_fd_sc_hd__a221o_1 _2705_ (.A1(_1062_),
    .A2(_1064_),
    .B1(_1068_),
    .B2(_1070_),
    .C1(_0797_),
    .X(_1071_));
 sky130_fd_sc_hd__mux4_1 _2706_ (.A0(\tms1x00.RAM[108][2] ),
    .A1(\tms1x00.RAM[109][2] ),
    .A2(\tms1x00.RAM[110][2] ),
    .A3(\tms1x00.RAM[111][2] ),
    .S0(_0939_),
    .S1(_0933_),
    .X(_1072_));
 sky130_fd_sc_hd__or2_1 _2707_ (.A(_0997_),
    .B(_1072_),
    .X(_1073_));
 sky130_fd_sc_hd__mux4_1 _2708_ (.A0(\tms1x00.RAM[104][2] ),
    .A1(\tms1x00.RAM[105][2] ),
    .A2(\tms1x00.RAM[106][2] ),
    .A3(\tms1x00.RAM[107][2] ),
    .S0(_0844_),
    .S1(_0946_),
    .X(_1074_));
 sky130_fd_sc_hd__o21a_1 _2709_ (.A1(_0802_),
    .A2(_1074_),
    .B1(_0800_),
    .X(_1075_));
 sky130_fd_sc_hd__mux4_1 _2710_ (.A0(\tms1x00.RAM[96][2] ),
    .A1(\tms1x00.RAM[97][2] ),
    .A2(\tms1x00.RAM[98][2] ),
    .A3(\tms1x00.RAM[99][2] ),
    .S0(_0932_),
    .S1(_0946_),
    .X(_1076_));
 sky130_fd_sc_hd__or2_1 _2711_ (.A(_0777_),
    .B(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__mux4_1 _2712_ (.A0(\tms1x00.RAM[100][2] ),
    .A1(\tms1x00.RAM[101][2] ),
    .A2(\tms1x00.RAM[102][2] ),
    .A3(\tms1x00.RAM[103][2] ),
    .S0(_0803_),
    .S1(_0804_),
    .X(_1078_));
 sky130_fd_sc_hd__o21a_1 _2713_ (.A1(_0816_),
    .A2(_1078_),
    .B1(_0766_),
    .X(_1079_));
 sky130_fd_sc_hd__a221o_1 _2714_ (.A1(_1073_),
    .A2(_1075_),
    .B1(_1077_),
    .B2(_1079_),
    .C1(_0039_),
    .X(_1080_));
 sky130_fd_sc_hd__a31o_1 _2715_ (.A1(_0040_),
    .A2(_1071_),
    .A3(_1080_),
    .B1(_0827_),
    .X(_1081_));
 sky130_fd_sc_hd__a31o_1 _2716_ (.A1(_0764_),
    .A2(_1046_),
    .A3(_1060_),
    .B1(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__mux4_1 _2717_ (.A0(\tms1x00.RAM[16][2] ),
    .A1(\tms1x00.RAM[17][2] ),
    .A2(\tms1x00.RAM[18][2] ),
    .A3(\tms1x00.RAM[19][2] ),
    .S0(_0807_),
    .S1(_0781_),
    .X(_1083_));
 sky130_fd_sc_hd__mux4_1 _2718_ (.A0(\tms1x00.RAM[20][2] ),
    .A1(\tms1x00.RAM[21][2] ),
    .A2(\tms1x00.RAM[22][2] ),
    .A3(\tms1x00.RAM[23][2] ),
    .S0(_0807_),
    .S1(_0781_),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_1 _2719_ (.A0(_1083_),
    .A1(_1084_),
    .S(_0865_),
    .X(_1085_));
 sky130_fd_sc_hd__mux2_1 _2720_ (.A0(\tms1x00.RAM[28][2] ),
    .A1(\tms1x00.RAM[29][2] ),
    .S(_1042_),
    .X(_1086_));
 sky130_fd_sc_hd__mux2_1 _2721_ (.A0(\tms1x00.RAM[30][2] ),
    .A1(\tms1x00.RAM[31][2] ),
    .S(_0994_),
    .X(_1087_));
 sky130_fd_sc_hd__a21o_1 _2722_ (.A1(_1037_),
    .A2(_1087_),
    .B1(_0828_),
    .X(_1088_));
 sky130_fd_sc_hd__a21o_1 _2723_ (.A1(_0857_),
    .A2(_1086_),
    .B1(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__mux4_1 _2724_ (.A0(\tms1x00.RAM[24][2] ),
    .A1(\tms1x00.RAM[25][2] ),
    .A2(\tms1x00.RAM[26][2] ),
    .A3(\tms1x00.RAM[27][2] ),
    .S0(_0858_),
    .S1(_0860_),
    .X(_1090_));
 sky130_fd_sc_hd__o21a_1 _2725_ (.A1(_1044_),
    .A2(_1090_),
    .B1(_0801_),
    .X(_1091_));
 sky130_fd_sc_hd__a221o_1 _2726_ (.A1(_0767_),
    .A2(_1085_),
    .B1(_1089_),
    .B2(_1091_),
    .C1(_0798_),
    .X(_1092_));
 sky130_fd_sc_hd__mux4_1 _2727_ (.A0(\tms1x00.RAM[8][2] ),
    .A1(\tms1x00.RAM[9][2] ),
    .A2(\tms1x00.RAM[10][2] ),
    .A3(\tms1x00.RAM[11][2] ),
    .S0(_1047_),
    .S1(_0938_),
    .X(_1093_));
 sky130_fd_sc_hd__or2_1 _2728_ (.A(_0865_),
    .B(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__or2b_1 _2729_ (.A(\tms1x00.RAM[15][2] ),
    .B_N(_1042_),
    .X(_1095_));
 sky130_fd_sc_hd__o21a_1 _2730_ (.A1(_1042_),
    .A2(\tms1x00.RAM[14][2] ),
    .B1(_1037_),
    .X(_1096_));
 sky130_fd_sc_hd__mux2_1 _2731_ (.A0(\tms1x00.RAM[12][2] ),
    .A1(\tms1x00.RAM[13][2] ),
    .S(_1042_),
    .X(_1097_));
 sky130_fd_sc_hd__a221o_1 _2732_ (.A1(_1095_),
    .A2(_1096_),
    .B1(_1097_),
    .B2(_0857_),
    .C1(_0828_),
    .X(_1098_));
 sky130_fd_sc_hd__mux2_1 _2733_ (.A0(\tms1x00.RAM[6][2] ),
    .A1(\tms1x00.RAM[7][2] ),
    .S(_0833_),
    .X(_1099_));
 sky130_fd_sc_hd__and2_1 _2734_ (.A(_1037_),
    .B(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_1 _2735_ (.A0(\tms1x00.RAM[4][2] ),
    .A1(\tms1x00.RAM[5][2] ),
    .S(_0812_),
    .X(_1101_));
 sky130_fd_sc_hd__a21o_1 _2736_ (.A1(_0814_),
    .A2(_1101_),
    .B1(_0997_),
    .X(_1102_));
 sky130_fd_sc_hd__mux4_1 _2737_ (.A0(\tms1x00.RAM[0][2] ),
    .A1(\tms1x00.RAM[1][2] ),
    .A2(\tms1x00.RAM[2][2] ),
    .A3(\tms1x00.RAM[3][2] ),
    .S0(_1047_),
    .S1(_0938_),
    .X(_1103_));
 sky130_fd_sc_hd__o221a_1 _2738_ (.A1(_1100_),
    .A2(_1102_),
    .B1(_1103_),
    .B2(_1044_),
    .C1(_0824_),
    .X(_1104_));
 sky130_fd_sc_hd__a311o_1 _2739_ (.A1(_0801_),
    .A2(_1094_),
    .A3(_1098_),
    .B1(_0818_),
    .C1(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__mux4_1 _2740_ (.A0(\tms1x00.RAM[44][2] ),
    .A1(\tms1x00.RAM[45][2] ),
    .A2(\tms1x00.RAM[46][2] ),
    .A3(\tms1x00.RAM[47][2] ),
    .S0(_0939_),
    .S1(_0780_),
    .X(_1106_));
 sky130_fd_sc_hd__or2_1 _2741_ (.A(_0862_),
    .B(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__mux4_1 _2742_ (.A0(\tms1x00.RAM[40][2] ),
    .A1(\tms1x00.RAM[41][2] ),
    .A2(\tms1x00.RAM[42][2] ),
    .A3(\tms1x00.RAM[43][2] ),
    .S0(_0932_),
    .S1(_0933_),
    .X(_1108_));
 sky130_fd_sc_hd__o21a_1 _2743_ (.A1(_0777_),
    .A2(_1108_),
    .B1(_0800_),
    .X(_1109_));
 sky130_fd_sc_hd__mux4_1 _2744_ (.A0(\tms1x00.RAM[32][2] ),
    .A1(\tms1x00.RAM[33][2] ),
    .A2(\tms1x00.RAM[34][2] ),
    .A3(\tms1x00.RAM[35][2] ),
    .S0(_0939_),
    .S1(_0933_),
    .X(_1110_));
 sky130_fd_sc_hd__or2_1 _2745_ (.A(_0777_),
    .B(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__mux4_2 _2746_ (.A0(\tms1x00.RAM[36][2] ),
    .A1(\tms1x00.RAM[37][2] ),
    .A2(\tms1x00.RAM[38][2] ),
    .A3(\tms1x00.RAM[39][2] ),
    .S0(_0932_),
    .S1(_0946_),
    .X(_1112_));
 sky130_fd_sc_hd__o21a_1 _2747_ (.A1(_0997_),
    .A2(_1112_),
    .B1(_0766_),
    .X(_1113_));
 sky130_fd_sc_hd__a221o_1 _2748_ (.A1(_1107_),
    .A2(_1109_),
    .B1(_1111_),
    .B2(_1113_),
    .C1(_0039_),
    .X(_1114_));
 sky130_fd_sc_hd__mux4_1 _2749_ (.A0(\tms1x00.RAM[56][2] ),
    .A1(\tms1x00.RAM[57][2] ),
    .A2(\tms1x00.RAM[58][2] ),
    .A3(\tms1x00.RAM[59][2] ),
    .S0(_0939_),
    .S1(_0780_),
    .X(_1115_));
 sky130_fd_sc_hd__or2_1 _2750_ (.A(_0777_),
    .B(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__mux4_1 _2751_ (.A0(\tms1x00.RAM[60][2] ),
    .A1(\tms1x00.RAM[61][2] ),
    .A2(\tms1x00.RAM[62][2] ),
    .A3(\tms1x00.RAM[63][2] ),
    .S0(_0932_),
    .S1(_0933_),
    .X(_1117_));
 sky130_fd_sc_hd__o21a_1 _2752_ (.A1(_0997_),
    .A2(_1117_),
    .B1(_0800_),
    .X(_1118_));
 sky130_fd_sc_hd__or2b_1 _2753_ (.A(\tms1x00.RAM[55][2] ),
    .B_N(_0994_),
    .X(_1119_));
 sky130_fd_sc_hd__o21a_1 _2754_ (.A1(_0873_),
    .A2(\tms1x00.RAM[54][2] ),
    .B1(_0771_),
    .X(_1120_));
 sky130_fd_sc_hd__mux2_1 _2755_ (.A0(\tms1x00.RAM[52][2] ),
    .A1(\tms1x00.RAM[53][2] ),
    .S(_0833_),
    .X(_1121_));
 sky130_fd_sc_hd__a221o_1 _2756_ (.A1(_1119_),
    .A2(_1120_),
    .B1(_1121_),
    .B2(_0814_),
    .C1(_0997_),
    .X(_1122_));
 sky130_fd_sc_hd__mux4_1 _2757_ (.A0(\tms1x00.RAM[48][2] ),
    .A1(\tms1x00.RAM[49][2] ),
    .A2(\tms1x00.RAM[50][2] ),
    .A3(\tms1x00.RAM[51][2] ),
    .S0(_0932_),
    .S1(_0946_),
    .X(_1123_));
 sky130_fd_sc_hd__o21a_1 _2758_ (.A1(_0802_),
    .A2(_1123_),
    .B1(_0766_),
    .X(_1124_));
 sky130_fd_sc_hd__a221o_1 _2759_ (.A1(_1116_),
    .A2(_1118_),
    .B1(_1122_),
    .B2(_1124_),
    .C1(_0797_),
    .X(_1125_));
 sky130_fd_sc_hd__a31o_1 _2760_ (.A1(_0040_),
    .A2(_1114_),
    .A3(_1125_),
    .B1(_0041_),
    .X(_1126_));
 sky130_fd_sc_hd__a31o_2 _2761_ (.A1(_0764_),
    .A2(_1092_),
    .A3(_1105_),
    .B1(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__a21oi_1 _2762_ (.A1(_1082_),
    .A2(_1127_),
    .B1(_0756_),
    .Y(_1128_));
 sky130_fd_sc_hd__a31o_1 _2763_ (.A1(_0742_),
    .A2(_0763_),
    .A3(_0909_),
    .B1(_0914_),
    .X(_1129_));
 sky130_fd_sc_hd__nand2_1 _2764_ (.A(\tms1x00.A[2] ),
    .B(_0931_),
    .Y(_1130_));
 sky130_fd_sc_hd__o21ai_4 _2765_ (.A1(_1128_),
    .A2(_1129_),
    .B1(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__buf_4 _2766_ (.A(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__buf_4 _2767_ (.A(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _2768_ (.A0(\tms1x00.RAM[109][2] ),
    .A1(_1133_),
    .S(_0929_),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _2769_ (.A(_1134_),
    .X(_0053_));
 sky130_fd_sc_hd__nand2_1 _2770_ (.A(_0742_),
    .B(\tms1x00.ins_in[6] ),
    .Y(_1135_));
 sky130_fd_sc_hd__inv_2 _2771_ (.A(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__mux4_1 _2772_ (.A0(\tms1x00.RAM[16][3] ),
    .A1(\tms1x00.RAM[17][3] ),
    .A2(\tms1x00.RAM[18][3] ),
    .A3(\tms1x00.RAM[19][3] ),
    .S0(_0858_),
    .S1(_0860_),
    .X(_1137_));
 sky130_fd_sc_hd__mux4_1 _2773_ (.A0(\tms1x00.RAM[20][3] ),
    .A1(\tms1x00.RAM[21][3] ),
    .A2(\tms1x00.RAM[22][3] ),
    .A3(\tms1x00.RAM[23][3] ),
    .S0(_1047_),
    .S1(_0860_),
    .X(_1138_));
 sky130_fd_sc_hd__mux2_1 _2774_ (.A0(_1137_),
    .A1(_1138_),
    .S(_0865_),
    .X(_1139_));
 sky130_fd_sc_hd__mux2_1 _2775_ (.A0(\tms1x00.RAM[30][3] ),
    .A1(\tms1x00.RAM[31][3] ),
    .S(_0812_),
    .X(_1140_));
 sky130_fd_sc_hd__and2_1 _2776_ (.A(_1037_),
    .B(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__mux2_1 _2777_ (.A0(\tms1x00.RAM[28][3] ),
    .A1(\tms1x00.RAM[29][3] ),
    .S(_0873_),
    .X(_1142_));
 sky130_fd_sc_hd__a21o_1 _2778_ (.A1(_0857_),
    .A2(_1142_),
    .B1(_0816_),
    .X(_1143_));
 sky130_fd_sc_hd__mux4_1 _2779_ (.A0(\tms1x00.RAM[24][3] ),
    .A1(\tms1x00.RAM[25][3] ),
    .A2(\tms1x00.RAM[26][3] ),
    .A3(\tms1x00.RAM[27][3] ),
    .S0(_0858_),
    .S1(_0860_),
    .X(_1144_));
 sky130_fd_sc_hd__o221a_1 _2780_ (.A1(_1141_),
    .A2(_1143_),
    .B1(_1144_),
    .B2(_1044_),
    .C1(_0801_),
    .X(_1145_));
 sky130_fd_sc_hd__a211o_1 _2781_ (.A1(_0767_),
    .A2(_1139_),
    .B1(_1145_),
    .C1(_0798_),
    .X(_1146_));
 sky130_fd_sc_hd__mux2_1 _2782_ (.A0(\tms1x00.RAM[6][3] ),
    .A1(\tms1x00.RAM[7][3] ),
    .S(_0774_),
    .X(_1147_));
 sky130_fd_sc_hd__and2_1 _2783_ (.A(_0860_),
    .B(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__mux2_1 _2784_ (.A0(\tms1x00.RAM[4][3] ),
    .A1(\tms1x00.RAM[5][3] ),
    .S(_0833_),
    .X(_1149_));
 sky130_fd_sc_hd__a21o_1 _2785_ (.A1(_0814_),
    .A2(_1149_),
    .B1(_0862_),
    .X(_1150_));
 sky130_fd_sc_hd__mux4_1 _2786_ (.A0(\tms1x00.RAM[0][3] ),
    .A1(\tms1x00.RAM[1][3] ),
    .A2(\tms1x00.RAM[2][3] ),
    .A3(\tms1x00.RAM[3][3] ),
    .S0(_0807_),
    .S1(_0781_),
    .X(_1151_));
 sky130_fd_sc_hd__o221a_1 _2787_ (.A1(_1148_),
    .A2(_1150_),
    .B1(_1151_),
    .B2(_0865_),
    .C1(_0824_),
    .X(_1152_));
 sky130_fd_sc_hd__mux4_1 _2788_ (.A0(\tms1x00.RAM[8][3] ),
    .A1(\tms1x00.RAM[9][3] ),
    .A2(\tms1x00.RAM[10][3] ),
    .A3(\tms1x00.RAM[11][3] ),
    .S0(_1047_),
    .S1(_0938_),
    .X(_1153_));
 sky130_fd_sc_hd__or2b_1 _2789_ (.A(\tms1x00.RAM[15][3] ),
    .B_N(_0873_),
    .X(_1154_));
 sky130_fd_sc_hd__o21a_1 _2790_ (.A1(_0873_),
    .A2(\tms1x00.RAM[14][3] ),
    .B1(_0804_),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _2791_ (.A0(\tms1x00.RAM[12][3] ),
    .A1(\tms1x00.RAM[13][3] ),
    .S(_0833_),
    .X(_1156_));
 sky130_fd_sc_hd__a221o_1 _2792_ (.A1(_1154_),
    .A2(_1155_),
    .B1(_1156_),
    .B2(_0814_),
    .C1(_0862_),
    .X(_1157_));
 sky130_fd_sc_hd__o211a_1 _2793_ (.A1(_1044_),
    .A2(_1153_),
    .B1(_1157_),
    .C1(_0795_),
    .X(_1158_));
 sky130_fd_sc_hd__or3_1 _2794_ (.A(_0818_),
    .B(_1152_),
    .C(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__mux4_1 _2795_ (.A0(\tms1x00.RAM[44][3] ),
    .A1(\tms1x00.RAM[45][3] ),
    .A2(\tms1x00.RAM[46][3] ),
    .A3(\tms1x00.RAM[47][3] ),
    .S0(_1047_),
    .S1(_0938_),
    .X(_1160_));
 sky130_fd_sc_hd__mux4_1 _2796_ (.A0(\tms1x00.RAM[40][3] ),
    .A1(\tms1x00.RAM[41][3] ),
    .A2(\tms1x00.RAM[42][3] ),
    .A3(\tms1x00.RAM[43][3] ),
    .S0(_0939_),
    .S1(_0933_),
    .X(_1161_));
 sky130_fd_sc_hd__or2_1 _2797_ (.A(_0777_),
    .B(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__o211a_1 _2798_ (.A1(_0828_),
    .A2(_1160_),
    .B1(_1162_),
    .C1(_0801_),
    .X(_1163_));
 sky130_fd_sc_hd__mux4_1 _2799_ (.A0(\tms1x00.RAM[32][3] ),
    .A1(\tms1x00.RAM[33][3] ),
    .A2(\tms1x00.RAM[34][3] ),
    .A3(\tms1x00.RAM[35][3] ),
    .S0(_1042_),
    .S1(_1037_),
    .X(_1164_));
 sky130_fd_sc_hd__mux4_1 _2800_ (.A0(\tms1x00.RAM[36][3] ),
    .A1(\tms1x00.RAM[37][3] ),
    .A2(\tms1x00.RAM[38][3] ),
    .A3(\tms1x00.RAM[39][3] ),
    .S0(_0844_),
    .S1(_0946_),
    .X(_1165_));
 sky130_fd_sc_hd__or2_1 _2801_ (.A(_0997_),
    .B(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__o211a_1 _2802_ (.A1(_1044_),
    .A2(_1164_),
    .B1(_1166_),
    .C1(_0767_),
    .X(_1167_));
 sky130_fd_sc_hd__mux4_1 _2803_ (.A0(\tms1x00.RAM[56][3] ),
    .A1(\tms1x00.RAM[57][3] ),
    .A2(\tms1x00.RAM[58][3] ),
    .A3(\tms1x00.RAM[59][3] ),
    .S0(_0803_),
    .S1(_0804_),
    .X(_1168_));
 sky130_fd_sc_hd__or2_1 _2804_ (.A(_0802_),
    .B(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__mux4_2 _2805_ (.A0(\tms1x00.RAM[60][3] ),
    .A1(\tms1x00.RAM[61][3] ),
    .A2(\tms1x00.RAM[62][3] ),
    .A3(\tms1x00.RAM[63][3] ),
    .S0(_0769_),
    .S1(_0771_),
    .X(_1170_));
 sky130_fd_sc_hd__o21a_1 _2806_ (.A1(_0828_),
    .A2(_1170_),
    .B1(_0800_),
    .X(_1171_));
 sky130_fd_sc_hd__or2b_1 _2807_ (.A(\tms1x00.RAM[55][3] ),
    .B_N(_1047_),
    .X(_1172_));
 sky130_fd_sc_hd__o21a_1 _2808_ (.A1(_1047_),
    .A2(\tms1x00.RAM[54][3] ),
    .B1(_0809_),
    .X(_1173_));
 sky130_fd_sc_hd__mux2_1 _2809_ (.A0(\tms1x00.RAM[52][3] ),
    .A1(\tms1x00.RAM[53][3] ),
    .S(_0873_),
    .X(_1174_));
 sky130_fd_sc_hd__a221o_1 _2810_ (.A1(_1172_),
    .A2(_1173_),
    .B1(_1174_),
    .B2(_0814_),
    .C1(_0816_),
    .X(_1175_));
 sky130_fd_sc_hd__mux4_2 _2811_ (.A0(\tms1x00.RAM[48][3] ),
    .A1(\tms1x00.RAM[49][3] ),
    .A2(\tms1x00.RAM[50][3] ),
    .A3(\tms1x00.RAM[51][3] ),
    .S0(_0769_),
    .S1(_0792_),
    .X(_1176_));
 sky130_fd_sc_hd__o21a_1 _2812_ (.A1(_0794_),
    .A2(_1176_),
    .B1(_0766_),
    .X(_1177_));
 sky130_fd_sc_hd__a221o_1 _2813_ (.A1(_1169_),
    .A2(_1171_),
    .B1(_1175_),
    .B2(_1177_),
    .C1(_0798_),
    .X(_1178_));
 sky130_fd_sc_hd__o311a_1 _2814_ (.A1(_0818_),
    .A2(_1163_),
    .A3(_1167_),
    .B1(_0040_),
    .C1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__a31o_1 _2815_ (.A1(_0764_),
    .A2(_1146_),
    .A3(_1159_),
    .B1(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__mux4_1 _2816_ (.A0(\tms1x00.RAM[80][3] ),
    .A1(\tms1x00.RAM[81][3] ),
    .A2(\tms1x00.RAM[82][3] ),
    .A3(\tms1x00.RAM[83][3] ),
    .S0(_0994_),
    .S1(_0781_),
    .X(_1181_));
 sky130_fd_sc_hd__mux4_1 _2817_ (.A0(\tms1x00.RAM[84][3] ),
    .A1(\tms1x00.RAM[85][3] ),
    .A2(\tms1x00.RAM[86][3] ),
    .A3(\tms1x00.RAM[87][3] ),
    .S0(_0994_),
    .S1(_0781_),
    .X(_1182_));
 sky130_fd_sc_hd__mux2_1 _2818_ (.A0(_1181_),
    .A1(_1182_),
    .S(_0865_),
    .X(_1183_));
 sky130_fd_sc_hd__mux2_1 _2819_ (.A0(\tms1x00.RAM[92][3] ),
    .A1(\tms1x00.RAM[93][3] ),
    .S(_1042_),
    .X(_1184_));
 sky130_fd_sc_hd__mux2_1 _2820_ (.A0(\tms1x00.RAM[94][3] ),
    .A1(\tms1x00.RAM[95][3] ),
    .S(_0994_),
    .X(_1185_));
 sky130_fd_sc_hd__a21o_1 _2821_ (.A1(_1037_),
    .A2(_1185_),
    .B1(_0828_),
    .X(_1186_));
 sky130_fd_sc_hd__a21o_1 _2822_ (.A1(_0857_),
    .A2(_1184_),
    .B1(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__mux4_1 _2823_ (.A0(\tms1x00.RAM[88][3] ),
    .A1(\tms1x00.RAM[89][3] ),
    .A2(\tms1x00.RAM[90][3] ),
    .A3(\tms1x00.RAM[91][3] ),
    .S0(_0858_),
    .S1(_0860_),
    .X(_1188_));
 sky130_fd_sc_hd__o21a_1 _2824_ (.A1(_1044_),
    .A2(_1188_),
    .B1(_0795_),
    .X(_1189_));
 sky130_fd_sc_hd__a221o_1 _2825_ (.A1(_0767_),
    .A2(_1183_),
    .B1(_1187_),
    .B2(_1189_),
    .C1(_0798_),
    .X(_1190_));
 sky130_fd_sc_hd__mux2_1 _2826_ (.A0(\tms1x00.RAM[70][3] ),
    .A1(\tms1x00.RAM[71][3] ),
    .S(_0844_),
    .X(_1191_));
 sky130_fd_sc_hd__and2_1 _2827_ (.A(_0938_),
    .B(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__mux2_1 _2828_ (.A0(\tms1x00.RAM[68][3] ),
    .A1(\tms1x00.RAM[69][3] ),
    .S(_0774_),
    .X(_1193_));
 sky130_fd_sc_hd__a21o_1 _2829_ (.A1(_0786_),
    .A2(_1193_),
    .B1(_0862_),
    .X(_1194_));
 sky130_fd_sc_hd__mux4_1 _2830_ (.A0(\tms1x00.RAM[64][3] ),
    .A1(\tms1x00.RAM[65][3] ),
    .A2(\tms1x00.RAM[66][3] ),
    .A3(\tms1x00.RAM[67][3] ),
    .S0(_0873_),
    .S1(_0781_),
    .X(_1195_));
 sky130_fd_sc_hd__o221a_1 _2831_ (.A1(_1192_),
    .A2(_1194_),
    .B1(_1195_),
    .B2(_0865_),
    .C1(_0824_),
    .X(_1196_));
 sky130_fd_sc_hd__mux4_1 _2832_ (.A0(\tms1x00.RAM[72][3] ),
    .A1(\tms1x00.RAM[73][3] ),
    .A2(\tms1x00.RAM[74][3] ),
    .A3(\tms1x00.RAM[75][3] ),
    .S0(_0807_),
    .S1(_0938_),
    .X(_1197_));
 sky130_fd_sc_hd__or2b_1 _2833_ (.A(\tms1x00.RAM[79][3] ),
    .B_N(_0873_),
    .X(_1198_));
 sky130_fd_sc_hd__o21a_1 _2834_ (.A1(_0873_),
    .A2(\tms1x00.RAM[78][3] ),
    .B1(_0946_),
    .X(_1199_));
 sky130_fd_sc_hd__mux2_1 _2835_ (.A0(\tms1x00.RAM[76][3] ),
    .A1(\tms1x00.RAM[77][3] ),
    .S(_0769_),
    .X(_1200_));
 sky130_fd_sc_hd__a221o_1 _2836_ (.A1(_1198_),
    .A2(_1199_),
    .B1(_1200_),
    .B2(_0786_),
    .C1(_0862_),
    .X(_1201_));
 sky130_fd_sc_hd__o211a_1 _2837_ (.A1(_0865_),
    .A2(_1197_),
    .B1(_1201_),
    .C1(_0795_),
    .X(_1202_));
 sky130_fd_sc_hd__or3_1 _2838_ (.A(_0818_),
    .B(_1196_),
    .C(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__mux4_1 _2839_ (.A0(\tms1x00.RAM[124][3] ),
    .A1(\tms1x00.RAM[125][3] ),
    .A2(\tms1x00.RAM[126][3] ),
    .A3(\tms1x00.RAM[127][3] ),
    .S0(_1047_),
    .S1(_0938_),
    .X(_1204_));
 sky130_fd_sc_hd__mux4_1 _2840_ (.A0(\tms1x00.RAM[120][3] ),
    .A1(\tms1x00.RAM[121][3] ),
    .A2(\tms1x00.RAM[122][3] ),
    .A3(\tms1x00.RAM[123][3] ),
    .S0(_0787_),
    .S1(_0780_),
    .X(_1205_));
 sky130_fd_sc_hd__or2_1 _2841_ (.A(_0848_),
    .B(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__o211a_1 _2842_ (.A1(_0828_),
    .A2(_1204_),
    .B1(_1206_),
    .C1(_0795_),
    .X(_1207_));
 sky130_fd_sc_hd__mux4_1 _2843_ (.A0(\tms1x00.RAM[112][3] ),
    .A1(\tms1x00.RAM[113][3] ),
    .A2(\tms1x00.RAM[114][3] ),
    .A3(\tms1x00.RAM[115][3] ),
    .S0(_1047_),
    .S1(_0938_),
    .X(_1208_));
 sky130_fd_sc_hd__or2b_1 _2844_ (.A(\tms1x00.RAM[119][3] ),
    .B_N(_0994_),
    .X(_1209_));
 sky130_fd_sc_hd__o21a_1 _2845_ (.A1(_0994_),
    .A2(\tms1x00.RAM[118][3] ),
    .B1(_0792_),
    .X(_1210_));
 sky130_fd_sc_hd__mux2_1 _2846_ (.A0(\tms1x00.RAM[116][3] ),
    .A1(\tms1x00.RAM[117][3] ),
    .S(_0833_),
    .X(_1211_));
 sky130_fd_sc_hd__a221o_1 _2847_ (.A1(_1209_),
    .A2(_1210_),
    .B1(_1211_),
    .B2(_0814_),
    .C1(_0997_),
    .X(_1212_));
 sky130_fd_sc_hd__o211a_1 _2848_ (.A1(_1044_),
    .A2(_1208_),
    .B1(_1212_),
    .C1(_0824_),
    .X(_1213_));
 sky130_fd_sc_hd__mux4_1 _2849_ (.A0(\tms1x00.RAM[108][3] ),
    .A1(\tms1x00.RAM[109][3] ),
    .A2(\tms1x00.RAM[110][3] ),
    .A3(\tms1x00.RAM[111][3] ),
    .S0(_0939_),
    .S1(_0933_),
    .X(_1214_));
 sky130_fd_sc_hd__or2_1 _2850_ (.A(_0997_),
    .B(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__mux4_1 _2851_ (.A0(\tms1x00.RAM[104][3] ),
    .A1(\tms1x00.RAM[105][3] ),
    .A2(\tms1x00.RAM[106][3] ),
    .A3(\tms1x00.RAM[107][3] ),
    .S0(_0844_),
    .S1(_0946_),
    .X(_1216_));
 sky130_fd_sc_hd__o21a_1 _2852_ (.A1(_0802_),
    .A2(_1216_),
    .B1(_0800_),
    .X(_1217_));
 sky130_fd_sc_hd__mux4_1 _2853_ (.A0(\tms1x00.RAM[96][3] ),
    .A1(\tms1x00.RAM[97][3] ),
    .A2(\tms1x00.RAM[98][3] ),
    .A3(\tms1x00.RAM[99][3] ),
    .S0(_0932_),
    .S1(_0933_),
    .X(_1218_));
 sky130_fd_sc_hd__or2_1 _2854_ (.A(_0777_),
    .B(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__mux4_1 _2855_ (.A0(\tms1x00.RAM[100][3] ),
    .A1(\tms1x00.RAM[101][3] ),
    .A2(\tms1x00.RAM[102][3] ),
    .A3(\tms1x00.RAM[103][3] ),
    .S0(_0803_),
    .S1(_0804_),
    .X(_1220_));
 sky130_fd_sc_hd__o21a_1 _2856_ (.A1(_0816_),
    .A2(_1220_),
    .B1(_0766_),
    .X(_1221_));
 sky130_fd_sc_hd__a221o_1 _2857_ (.A1(_1215_),
    .A2(_1217_),
    .B1(_1219_),
    .B2(_1221_),
    .C1(_0039_),
    .X(_1222_));
 sky130_fd_sc_hd__o311a_1 _2858_ (.A1(_0798_),
    .A2(_1207_),
    .A3(_1213_),
    .B1(_1222_),
    .C1(_0040_),
    .X(_1223_));
 sky130_fd_sc_hd__a311o_1 _2859_ (.A1(_0764_),
    .A2(_1190_),
    .A3(_1203_),
    .B1(_1223_),
    .C1(_0827_),
    .X(_1224_));
 sky130_fd_sc_hd__o21ai_4 _2860_ (.A1(_0041_),
    .A2(_1180_),
    .B1(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__a2bb2o_1 _2861_ (.A1_N(_1135_),
    .A2_N(_0909_),
    .B1(_0931_),
    .B2(\tms1x00.A[3] ),
    .X(_1226_));
 sky130_fd_sc_hd__o21bai_2 _2862_ (.A1(_1136_),
    .A2(_1225_),
    .B1_N(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__buf_4 _2863_ (.A(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__buf_4 _2864_ (.A(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__mux2_1 _2865_ (.A0(\tms1x00.RAM[109][3] ),
    .A1(_1229_),
    .S(_0929_),
    .X(_1230_));
 sky130_fd_sc_hd__clkbuf_1 _2866_ (.A(_1230_),
    .X(_0054_));
 sky130_fd_sc_hd__nand2_1 _2867_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[1] ),
    .Y(_1231_));
 sky130_fd_sc_hd__or4_1 _2868_ (.A(_0730_),
    .B(_0734_),
    .C(_0926_),
    .D(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__buf_4 _2869_ (.A(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__nor2_2 _2870_ (.A(_0922_),
    .B(_1233_),
    .Y(_1234_));
 sky130_fd_sc_hd__mux2_1 _2871_ (.A0(\tms1x00.RAM[99][0] ),
    .A1(_0920_),
    .S(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__clkbuf_1 _2872_ (.A(_1235_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2873_ (.A0(\tms1x00.RAM[99][1] ),
    .A1(_1032_),
    .S(_1234_),
    .X(_1236_));
 sky130_fd_sc_hd__clkbuf_1 _2874_ (.A(_1236_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2875_ (.A0(\tms1x00.RAM[99][2] ),
    .A1(_1133_),
    .S(_1234_),
    .X(_1237_));
 sky130_fd_sc_hd__clkbuf_1 _2876_ (.A(_1237_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2877_ (.A0(\tms1x00.RAM[99][3] ),
    .A1(_1229_),
    .S(_1234_),
    .X(_1238_));
 sky130_fd_sc_hd__clkbuf_1 _2878_ (.A(_1238_),
    .X(_0058_));
 sky130_fd_sc_hd__buf_4 _2879_ (.A(_0919_),
    .X(_1239_));
 sky130_fd_sc_hd__or3b_4 _2880_ (.A(\tms1x00.ram_addr_buff[5] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C_N(\tms1x00.ram_addr_buff[4] ),
    .X(_1240_));
 sky130_fd_sc_hd__buf_4 _2881_ (.A(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__nor2_4 _2882_ (.A(_0908_),
    .B(_0916_),
    .Y(_1242_));
 sky130_fd_sc_hd__or4_4 _2883_ (.A(_0730_),
    .B(_0734_),
    .C(_0923_),
    .D(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__or2_2 _2884_ (.A(_1241_),
    .B(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_1 _2885_ (.A0(_1239_),
    .A1(\tms1x00.RAM[17][0] ),
    .S(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__clkbuf_1 _2886_ (.A(_1245_),
    .X(_0059_));
 sky130_fd_sc_hd__buf_4 _2887_ (.A(_1031_),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_1 _2888_ (.A0(_1246_),
    .A1(\tms1x00.RAM[17][1] ),
    .S(_1244_),
    .X(_1247_));
 sky130_fd_sc_hd__clkbuf_1 _2889_ (.A(_1247_),
    .X(_0060_));
 sky130_fd_sc_hd__clkbuf_4 _2890_ (.A(_1132_),
    .X(_1248_));
 sky130_fd_sc_hd__mux2_1 _2891_ (.A0(_1248_),
    .A1(\tms1x00.RAM[17][2] ),
    .S(_1244_),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_1 _2892_ (.A(_1249_),
    .X(_0061_));
 sky130_fd_sc_hd__buf_4 _2893_ (.A(_1228_),
    .X(_1250_));
 sky130_fd_sc_hd__mux2_1 _2894_ (.A0(_1250_),
    .A1(\tms1x00.RAM[17][3] ),
    .S(_1244_),
    .X(_1251_));
 sky130_fd_sc_hd__clkbuf_1 _2895_ (.A(_1251_),
    .X(_0062_));
 sky130_fd_sc_hd__nand3b_4 _2896_ (.A_N(\tms1x00.ram_addr_buff[5] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C(\tms1x00.ram_addr_buff[4] ),
    .Y(_1252_));
 sky130_fd_sc_hd__buf_4 _2897_ (.A(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__or3b_1 _2898_ (.A(_0730_),
    .B(_1242_),
    .C_N(_0734_),
    .X(_1254_));
 sky130_fd_sc_hd__or2_4 _2899_ (.A(_0923_),
    .B(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__or2_2 _2900_ (.A(_1253_),
    .B(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__mux2_1 _2901_ (.A0(_1239_),
    .A1(\tms1x00.RAM[89][0] ),
    .S(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__clkbuf_1 _2902_ (.A(_1257_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _2903_ (.A0(_1246_),
    .A1(\tms1x00.RAM[89][1] ),
    .S(_1256_),
    .X(_1258_));
 sky130_fd_sc_hd__clkbuf_1 _2904_ (.A(_1258_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _2905_ (.A0(_1248_),
    .A1(\tms1x00.RAM[89][2] ),
    .S(_1256_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_1 _2906_ (.A(_1259_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _2907_ (.A0(_1250_),
    .A1(\tms1x00.RAM[89][3] ),
    .S(_1256_),
    .X(_1260_));
 sky130_fd_sc_hd__clkbuf_1 _2908_ (.A(_1260_),
    .X(_0066_));
 sky130_fd_sc_hd__or2_4 _2909_ (.A(_0924_),
    .B(_1231_),
    .X(_1261_));
 sky130_fd_sc_hd__or3b_1 _2910_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C_N(\tms1x00.ram_addr_buff[6] ),
    .X(_1262_));
 sky130_fd_sc_hd__buf_2 _2911_ (.A(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__or2_2 _2912_ (.A(_1242_),
    .B(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__or2_2 _2913_ (.A(_1261_),
    .B(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__mux2_1 _2914_ (.A0(_1239_),
    .A1(\tms1x00.RAM[79][0] ),
    .S(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__clkbuf_1 _2915_ (.A(_1266_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _2916_ (.A0(_1246_),
    .A1(\tms1x00.RAM[79][1] ),
    .S(_1265_),
    .X(_1267_));
 sky130_fd_sc_hd__clkbuf_1 _2917_ (.A(_1267_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2918_ (.A0(_1248_),
    .A1(\tms1x00.RAM[79][2] ),
    .S(_1265_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_1 _2919_ (.A(_1268_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _2920_ (.A0(_1250_),
    .A1(\tms1x00.RAM[79][3] ),
    .S(_1265_),
    .X(_1269_));
 sky130_fd_sc_hd__clkbuf_1 _2921_ (.A(_1269_),
    .X(_0070_));
 sky130_fd_sc_hd__or4b_1 _2922_ (.A(_0720_),
    .B(_0730_),
    .C(_0734_),
    .D_N(_0727_),
    .X(_1270_));
 sky130_fd_sc_hd__or2_4 _2923_ (.A(_1242_),
    .B(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__or2_2 _2924_ (.A(_1241_),
    .B(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__mux2_1 _2925_ (.A0(_1239_),
    .A1(\tms1x00.RAM[18][0] ),
    .S(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__clkbuf_1 _2926_ (.A(_1273_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _2927_ (.A0(_1246_),
    .A1(\tms1x00.RAM[18][1] ),
    .S(_1272_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _2928_ (.A(_1274_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _2929_ (.A0(_1248_),
    .A1(\tms1x00.RAM[18][2] ),
    .S(_1272_),
    .X(_1275_));
 sky130_fd_sc_hd__clkbuf_1 _2930_ (.A(_1275_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2931_ (.A0(_1250_),
    .A1(\tms1x00.RAM[18][3] ),
    .S(_1272_),
    .X(_1276_));
 sky130_fd_sc_hd__clkbuf_1 _2932_ (.A(_1276_),
    .X(_0074_));
 sky130_fd_sc_hd__or2b_1 _2933_ (.A(\tms1x00.ram_addr_buff[3] ),
    .B_N(\tms1x00.ram_addr_buff[2] ),
    .X(_1277_));
 sky130_fd_sc_hd__or3_4 _2934_ (.A(_0923_),
    .B(_1242_),
    .C(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__or2_2 _2935_ (.A(_1263_),
    .B(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__mux2_1 _2936_ (.A0(_1239_),
    .A1(\tms1x00.RAM[69][0] ),
    .S(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _2937_ (.A(_1280_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _2938_ (.A0(_1246_),
    .A1(\tms1x00.RAM[69][1] ),
    .S(_1279_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_1 _2939_ (.A(_1281_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2940_ (.A0(_1248_),
    .A1(\tms1x00.RAM[69][2] ),
    .S(_1279_),
    .X(_1282_));
 sky130_fd_sc_hd__clkbuf_1 _2941_ (.A(_1282_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2942_ (.A0(_1250_),
    .A1(\tms1x00.RAM[69][3] ),
    .S(_1279_),
    .X(_1283_));
 sky130_fd_sc_hd__clkbuf_1 _2943_ (.A(_1283_),
    .X(_0078_));
 sky130_fd_sc_hd__nand3b_2 _2944_ (.A_N(\tms1x00.ram_addr_buff[6] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[4] ),
    .Y(_1284_));
 sky130_fd_sc_hd__clkbuf_4 _2945_ (.A(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__clkbuf_4 _2946_ (.A(_0926_),
    .X(_1286_));
 sky130_fd_sc_hd__or3b_4 _2947_ (.A(_1231_),
    .B(_0730_),
    .C_N(_0734_),
    .X(_1287_));
 sky130_fd_sc_hd__or2_4 _2948_ (.A(_1286_),
    .B(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__or2_2 _2949_ (.A(_1285_),
    .B(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__mux2_1 _2950_ (.A0(_1239_),
    .A1(\tms1x00.RAM[59][0] ),
    .S(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _2951_ (.A(_1290_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _2952_ (.A0(_1246_),
    .A1(\tms1x00.RAM[59][1] ),
    .S(_1289_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _2953_ (.A(_1291_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2954_ (.A0(_1248_),
    .A1(\tms1x00.RAM[59][2] ),
    .S(_1289_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _2955_ (.A(_1292_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2956_ (.A0(_1250_),
    .A1(\tms1x00.RAM[59][3] ),
    .S(_1289_),
    .X(_1293_));
 sky130_fd_sc_hd__clkbuf_1 _2957_ (.A(_1293_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2958_ (.A0(\K_override[0] ),
    .A1(net68),
    .S(_0716_),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _2959_ (.A(_1294_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2960_ (.A0(\K_override[1] ),
    .A1(net69),
    .S(_0716_),
    .X(_1295_));
 sky130_fd_sc_hd__clkbuf_1 _2961_ (.A(_1295_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2962_ (.A0(\K_override[2] ),
    .A1(net63),
    .S(_0716_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _2963_ (.A(_1296_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2964_ (.A0(\K_override[3] ),
    .A1(net64),
    .S(_0716_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_1 _2965_ (.A(_1297_),
    .X(_0086_));
 sky130_fd_sc_hd__or2_2 _2966_ (.A(_1243_),
    .B(_1284_),
    .X(_1298_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(_1239_),
    .A1(\tms1x00.RAM[49][0] ),
    .S(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__clkbuf_1 _2968_ (.A(_1299_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2969_ (.A0(_1246_),
    .A1(\tms1x00.RAM[49][1] ),
    .S(_1298_),
    .X(_1300_));
 sky130_fd_sc_hd__clkbuf_1 _2970_ (.A(_1300_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2971_ (.A0(_1248_),
    .A1(\tms1x00.RAM[49][2] ),
    .S(_1298_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_1 _2972_ (.A(_1301_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2973_ (.A0(_1250_),
    .A1(\tms1x00.RAM[49][3] ),
    .S(_1298_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _2974_ (.A(_1302_),
    .X(_0090_));
 sky130_fd_sc_hd__nor2_2 _2975_ (.A(_1233_),
    .B(_1241_),
    .Y(_1303_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(\tms1x00.RAM[19][0] ),
    .A1(_0920_),
    .S(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_1 _2977_ (.A(_1304_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(\tms1x00.RAM[19][1] ),
    .A1(_1032_),
    .S(_1303_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_1 _2979_ (.A(_1305_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(\tms1x00.RAM[19][2] ),
    .A1(_1133_),
    .S(_1303_),
    .X(_1306_));
 sky130_fd_sc_hd__clkbuf_1 _2981_ (.A(_1306_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(\tms1x00.RAM[19][3] ),
    .A1(_1229_),
    .S(_1303_),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_1 _2983_ (.A(_1307_),
    .X(_0094_));
 sky130_fd_sc_hd__or4b_2 _2984_ (.A(_0720_),
    .B(_0727_),
    .C(_0730_),
    .D_N(_0734_),
    .X(_1308_));
 sky130_fd_sc_hd__or2_4 _2985_ (.A(_1286_),
    .B(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__nor2_2 _2986_ (.A(_0922_),
    .B(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__mux2_1 _2987_ (.A0(\tms1x00.RAM[104][0] ),
    .A1(_0920_),
    .S(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__clkbuf_1 _2988_ (.A(_1311_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(\tms1x00.RAM[104][1] ),
    .A1(_1032_),
    .S(_1310_),
    .X(_1312_));
 sky130_fd_sc_hd__clkbuf_1 _2990_ (.A(_1312_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _2991_ (.A0(\tms1x00.RAM[104][2] ),
    .A1(_1133_),
    .S(_1310_),
    .X(_1313_));
 sky130_fd_sc_hd__clkbuf_1 _2992_ (.A(_1313_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _2993_ (.A0(\tms1x00.RAM[104][3] ),
    .A1(_1229_),
    .S(_1310_),
    .X(_1314_));
 sky130_fd_sc_hd__clkbuf_1 _2994_ (.A(_1314_),
    .X(_0098_));
 sky130_fd_sc_hd__or2_1 _2995_ (.A(_1231_),
    .B(_1277_),
    .X(_1315_));
 sky130_fd_sc_hd__clkbuf_4 _2996_ (.A(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__nor3_2 _2997_ (.A(_0922_),
    .B(_1286_),
    .C(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__mux2_1 _2998_ (.A0(\tms1x00.RAM[103][0] ),
    .A1(_0920_),
    .S(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__clkbuf_1 _2999_ (.A(_1318_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _3000_ (.A0(\tms1x00.RAM[103][1] ),
    .A1(_1032_),
    .S(_1317_),
    .X(_1319_));
 sky130_fd_sc_hd__clkbuf_1 _3001_ (.A(_1319_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _3002_ (.A0(\tms1x00.RAM[103][2] ),
    .A1(_1133_),
    .S(_1317_),
    .X(_1320_));
 sky130_fd_sc_hd__clkbuf_1 _3003_ (.A(_1320_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _3004_ (.A0(\tms1x00.RAM[103][3] ),
    .A1(_1229_),
    .S(_1317_),
    .X(_1321_));
 sky130_fd_sc_hd__clkbuf_1 _3005_ (.A(_1321_),
    .X(_0102_));
 sky130_fd_sc_hd__or3b_2 _3006_ (.A(_1277_),
    .B(_0720_),
    .C_N(_0727_),
    .X(_1322_));
 sky130_fd_sc_hd__or2_1 _3007_ (.A(_1286_),
    .B(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__buf_6 _3008_ (.A(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__nor2_2 _3009_ (.A(_0922_),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__mux2_1 _3010_ (.A0(\tms1x00.RAM[102][0] ),
    .A1(_0920_),
    .S(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__clkbuf_1 _3011_ (.A(_1326_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _3012_ (.A0(\tms1x00.RAM[102][1] ),
    .A1(_1032_),
    .S(_1325_),
    .X(_1327_));
 sky130_fd_sc_hd__clkbuf_1 _3013_ (.A(_1327_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _3014_ (.A0(\tms1x00.RAM[102][2] ),
    .A1(_1133_),
    .S(_1325_),
    .X(_1328_));
 sky130_fd_sc_hd__clkbuf_1 _3015_ (.A(_1328_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _3016_ (.A0(\tms1x00.RAM[102][3] ),
    .A1(_1229_),
    .S(_1325_),
    .X(_1329_));
 sky130_fd_sc_hd__clkbuf_1 _3017_ (.A(_1329_),
    .X(_0106_));
 sky130_fd_sc_hd__or2_2 _3018_ (.A(_0922_),
    .B(_1278_),
    .X(_1330_));
 sky130_fd_sc_hd__mux2_1 _3019_ (.A0(_1239_),
    .A1(\tms1x00.RAM[101][0] ),
    .S(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__clkbuf_1 _3020_ (.A(_1331_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _3021_ (.A0(_1246_),
    .A1(\tms1x00.RAM[101][1] ),
    .S(_1330_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_1 _3022_ (.A(_1332_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _3023_ (.A0(_1248_),
    .A1(\tms1x00.RAM[101][2] ),
    .S(_1330_),
    .X(_1333_));
 sky130_fd_sc_hd__clkbuf_1 _3024_ (.A(_1333_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _3025_ (.A0(_1250_),
    .A1(\tms1x00.RAM[101][3] ),
    .S(_1330_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_1 _3026_ (.A(_1334_),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_8 _3027_ (.A(_0918_),
    .X(_1335_));
 sky130_fd_sc_hd__buf_4 _3028_ (.A(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__or3_2 _3029_ (.A(_0720_),
    .B(_0727_),
    .C(_1277_),
    .X(_1337_));
 sky130_fd_sc_hd__or2_1 _3030_ (.A(_1286_),
    .B(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__buf_4 _3031_ (.A(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__nor2_2 _3032_ (.A(_0922_),
    .B(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__mux2_1 _3033_ (.A0(\tms1x00.RAM[100][0] ),
    .A1(_1336_),
    .S(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__clkbuf_1 _3034_ (.A(_1341_),
    .X(_0111_));
 sky130_fd_sc_hd__buf_4 _3035_ (.A(_1030_),
    .X(_1342_));
 sky130_fd_sc_hd__buf_4 _3036_ (.A(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__mux2_1 _3037_ (.A0(\tms1x00.RAM[100][1] ),
    .A1(_1343_),
    .S(_1340_),
    .X(_1344_));
 sky130_fd_sc_hd__clkbuf_1 _3038_ (.A(_1344_),
    .X(_0112_));
 sky130_fd_sc_hd__buf_4 _3039_ (.A(_1131_),
    .X(_1345_));
 sky130_fd_sc_hd__buf_4 _3040_ (.A(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__mux2_1 _3041_ (.A0(\tms1x00.RAM[100][2] ),
    .A1(_1346_),
    .S(_1340_),
    .X(_1347_));
 sky130_fd_sc_hd__clkbuf_1 _3042_ (.A(_1347_),
    .X(_0113_));
 sky130_fd_sc_hd__buf_4 _3043_ (.A(_1227_),
    .X(_1348_));
 sky130_fd_sc_hd__buf_4 _3044_ (.A(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__mux2_1 _3045_ (.A0(\tms1x00.RAM[100][3] ),
    .A1(_1349_),
    .S(_1340_),
    .X(_1350_));
 sky130_fd_sc_hd__clkbuf_1 _3046_ (.A(_1350_),
    .X(_0114_));
 sky130_fd_sc_hd__or3_1 _3047_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[6] ),
    .X(_1351_));
 sky130_fd_sc_hd__clkbuf_4 _3048_ (.A(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__or4_4 _3049_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[1] ),
    .C(\tms1x00.ram_addr_buff[2] ),
    .D(\tms1x00.ram_addr_buff[3] ),
    .X(_1353_));
 sky130_fd_sc_hd__or2_1 _3050_ (.A(_1286_),
    .B(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__buf_4 _3051_ (.A(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__nor2_2 _3052_ (.A(_1352_),
    .B(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__mux2_1 _3053_ (.A0(\tms1x00.RAM[0][0] ),
    .A1(_1336_),
    .S(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__clkbuf_1 _3054_ (.A(_1357_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _3055_ (.A0(\tms1x00.RAM[0][1] ),
    .A1(_1343_),
    .S(_1356_),
    .X(_1358_));
 sky130_fd_sc_hd__clkbuf_1 _3056_ (.A(_1358_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _3057_ (.A0(\tms1x00.RAM[0][2] ),
    .A1(_1346_),
    .S(_1356_),
    .X(_1359_));
 sky130_fd_sc_hd__clkbuf_1 _3058_ (.A(_1359_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(\tms1x00.RAM[0][3] ),
    .A1(_1349_),
    .S(_1356_),
    .X(_1360_));
 sky130_fd_sc_hd__clkbuf_1 _3060_ (.A(_1360_),
    .X(_0118_));
 sky130_fd_sc_hd__or2_2 _3061_ (.A(_0922_),
    .B(_1271_),
    .X(_1361_));
 sky130_fd_sc_hd__mux2_1 _3062_ (.A0(_1239_),
    .A1(\tms1x00.RAM[98][0] ),
    .S(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _3063_ (.A(_1362_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _3064_ (.A0(_1246_),
    .A1(\tms1x00.RAM[98][1] ),
    .S(_1361_),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_1 _3065_ (.A(_1363_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _3066_ (.A0(_1248_),
    .A1(\tms1x00.RAM[98][2] ),
    .S(_1361_),
    .X(_1364_));
 sky130_fd_sc_hd__clkbuf_1 _3067_ (.A(_1364_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _3068_ (.A0(_1250_),
    .A1(\tms1x00.RAM[98][3] ),
    .S(_1361_),
    .X(_1365_));
 sky130_fd_sc_hd__clkbuf_1 _3069_ (.A(_1365_),
    .X(_0122_));
 sky130_fd_sc_hd__or2_2 _3070_ (.A(_0922_),
    .B(_1243_),
    .X(_1366_));
 sky130_fd_sc_hd__mux2_1 _3071_ (.A0(_1239_),
    .A1(\tms1x00.RAM[97][0] ),
    .S(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__clkbuf_1 _3072_ (.A(_1367_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _3073_ (.A0(_1246_),
    .A1(\tms1x00.RAM[97][1] ),
    .S(_1366_),
    .X(_1368_));
 sky130_fd_sc_hd__clkbuf_1 _3074_ (.A(_1368_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _3075_ (.A0(_1248_),
    .A1(\tms1x00.RAM[97][2] ),
    .S(_1366_),
    .X(_1369_));
 sky130_fd_sc_hd__clkbuf_1 _3076_ (.A(_1369_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _3077_ (.A0(_1250_),
    .A1(\tms1x00.RAM[97][3] ),
    .S(_1366_),
    .X(_1370_));
 sky130_fd_sc_hd__clkbuf_1 _3078_ (.A(_1370_),
    .X(_0126_));
 sky130_fd_sc_hd__nor2_2 _3079_ (.A(_0922_),
    .B(_1355_),
    .Y(_1371_));
 sky130_fd_sc_hd__mux2_1 _3080_ (.A0(\tms1x00.RAM[96][0] ),
    .A1(_1336_),
    .S(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__clkbuf_1 _3081_ (.A(_1372_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _3082_ (.A0(\tms1x00.RAM[96][1] ),
    .A1(_1343_),
    .S(_1371_),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_1 _3083_ (.A(_1373_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _3084_ (.A0(\tms1x00.RAM[96][2] ),
    .A1(_1346_),
    .S(_1371_),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_1 _3085_ (.A(_1374_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _3086_ (.A0(\tms1x00.RAM[96][3] ),
    .A1(_1349_),
    .S(_1371_),
    .X(_1375_));
 sky130_fd_sc_hd__clkbuf_1 _3087_ (.A(_1375_),
    .X(_0130_));
 sky130_fd_sc_hd__nor3_4 _3088_ (.A(_1242_),
    .B(_1253_),
    .C(_1261_),
    .Y(_1376_));
 sky130_fd_sc_hd__mux2_1 _3089_ (.A0(\tms1x00.RAM[95][0] ),
    .A1(_1336_),
    .S(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_1 _3090_ (.A(_1377_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _3091_ (.A0(\tms1x00.RAM[95][1] ),
    .A1(_1343_),
    .S(_1376_),
    .X(_1378_));
 sky130_fd_sc_hd__clkbuf_1 _3092_ (.A(_1378_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _3093_ (.A0(\tms1x00.RAM[95][2] ),
    .A1(_1346_),
    .S(_1376_),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _3094_ (.A(_1379_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _3095_ (.A0(\tms1x00.RAM[95][3] ),
    .A1(_1349_),
    .S(_1376_),
    .X(_1380_));
 sky130_fd_sc_hd__clkbuf_1 _3096_ (.A(_1380_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_4 _3097_ (.A(_0919_),
    .X(_1381_));
 sky130_fd_sc_hd__nand3_2 _3098_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[6] ),
    .Y(_1382_));
 sky130_fd_sc_hd__clkbuf_4 _3099_ (.A(_1382_),
    .X(_1383_));
 sky130_fd_sc_hd__or2_2 _3100_ (.A(_1271_),
    .B(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(_1381_),
    .A1(\tms1x00.RAM[114][0] ),
    .S(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__clkbuf_1 _3102_ (.A(_1385_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_4 _3103_ (.A(_1031_),
    .X(_1386_));
 sky130_fd_sc_hd__mux2_1 _3104_ (.A0(_1386_),
    .A1(\tms1x00.RAM[114][1] ),
    .S(_1384_),
    .X(_1387_));
 sky130_fd_sc_hd__clkbuf_1 _3105_ (.A(_1387_),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_4 _3106_ (.A(_1132_),
    .X(_1388_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(_1388_),
    .A1(\tms1x00.RAM[114][2] ),
    .S(_1384_),
    .X(_1389_));
 sky130_fd_sc_hd__clkbuf_1 _3108_ (.A(_1389_),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_4 _3109_ (.A(_1228_),
    .X(_1390_));
 sky130_fd_sc_hd__mux2_1 _3110_ (.A0(_1390_),
    .A1(\tms1x00.RAM[114][3] ),
    .S(_1384_),
    .X(_1391_));
 sky130_fd_sc_hd__clkbuf_1 _3111_ (.A(_1391_),
    .X(_0138_));
 sky130_fd_sc_hd__or2_2 _3112_ (.A(_1243_),
    .B(_1383_),
    .X(_1392_));
 sky130_fd_sc_hd__mux2_1 _3113_ (.A0(_1381_),
    .A1(\tms1x00.RAM[113][0] ),
    .S(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _3114_ (.A(_1393_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _3115_ (.A0(_1386_),
    .A1(\tms1x00.RAM[113][1] ),
    .S(_1392_),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _3116_ (.A(_1394_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _3117_ (.A0(_1388_),
    .A1(\tms1x00.RAM[113][2] ),
    .S(_1392_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_1 _3118_ (.A(_1395_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _3119_ (.A0(_1390_),
    .A1(\tms1x00.RAM[113][3] ),
    .S(_1392_),
    .X(_1396_));
 sky130_fd_sc_hd__clkbuf_1 _3120_ (.A(_1396_),
    .X(_0142_));
 sky130_fd_sc_hd__or2_2 _3121_ (.A(_1286_),
    .B(_1382_),
    .X(_1397_));
 sky130_fd_sc_hd__nor2_2 _3122_ (.A(_1353_),
    .B(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__mux2_1 _3123_ (.A0(\tms1x00.RAM[112][0] ),
    .A1(_1336_),
    .S(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_1 _3124_ (.A(_1399_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _3125_ (.A0(\tms1x00.RAM[112][1] ),
    .A1(_1343_),
    .S(_1398_),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_1 _3126_ (.A(_1400_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _3127_ (.A0(\tms1x00.RAM[112][2] ),
    .A1(_1346_),
    .S(_1398_),
    .X(_1401_));
 sky130_fd_sc_hd__clkbuf_1 _3128_ (.A(_1401_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _3129_ (.A0(\tms1x00.RAM[112][3] ),
    .A1(_1349_),
    .S(_1398_),
    .X(_1402_));
 sky130_fd_sc_hd__clkbuf_1 _3130_ (.A(_1402_),
    .X(_0146_));
 sky130_fd_sc_hd__or2_4 _3131_ (.A(_1286_),
    .B(_1261_),
    .X(_1403_));
 sky130_fd_sc_hd__or2_2 _3132_ (.A(_0921_),
    .B(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__mux2_1 _3133_ (.A0(_1381_),
    .A1(\tms1x00.RAM[111][0] ),
    .S(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_1 _3134_ (.A(_1405_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _3135_ (.A0(_1386_),
    .A1(\tms1x00.RAM[111][1] ),
    .S(_1404_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _3136_ (.A(_1406_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _3137_ (.A0(_1388_),
    .A1(\tms1x00.RAM[111][2] ),
    .S(_1404_),
    .X(_1407_));
 sky130_fd_sc_hd__clkbuf_1 _3138_ (.A(_1407_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _3139_ (.A0(_1390_),
    .A1(\tms1x00.RAM[111][3] ),
    .S(_1404_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _3140_ (.A(_1408_),
    .X(_0150_));
 sky130_fd_sc_hd__or2_1 _3141_ (.A(_0924_),
    .B(_1242_),
    .X(_1409_));
 sky130_fd_sc_hd__or3b_4 _3142_ (.A(_1409_),
    .B(_0720_),
    .C_N(_0727_),
    .X(_1410_));
 sky130_fd_sc_hd__or2_2 _3143_ (.A(_0921_),
    .B(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__mux2_1 _3144_ (.A0(_1381_),
    .A1(\tms1x00.RAM[110][0] ),
    .S(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__clkbuf_1 _3145_ (.A(_1412_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _3146_ (.A0(_1386_),
    .A1(\tms1x00.RAM[110][1] ),
    .S(_1411_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_1 _3147_ (.A(_1413_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _3148_ (.A0(_1388_),
    .A1(\tms1x00.RAM[110][2] ),
    .S(_1411_),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _3149_ (.A(_1414_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _3150_ (.A0(_1390_),
    .A1(\tms1x00.RAM[110][3] ),
    .S(_1411_),
    .X(_1415_));
 sky130_fd_sc_hd__clkbuf_1 _3151_ (.A(_1415_),
    .X(_0154_));
 sky130_fd_sc_hd__or3b_4 _3152_ (.A(_1254_),
    .B(_0720_),
    .C_N(_0727_),
    .X(_1416_));
 sky130_fd_sc_hd__or2_2 _3153_ (.A(_1352_),
    .B(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__mux2_1 _3154_ (.A0(_1381_),
    .A1(\tms1x00.RAM[10][0] ),
    .S(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _3155_ (.A(_1418_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _3156_ (.A0(_1386_),
    .A1(\tms1x00.RAM[10][1] ),
    .S(_1417_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_1 _3157_ (.A(_1419_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _3158_ (.A0(_1388_),
    .A1(\tms1x00.RAM[10][2] ),
    .S(_1417_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _3159_ (.A(_1420_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _3160_ (.A0(_1390_),
    .A1(\tms1x00.RAM[10][3] ),
    .S(_1417_),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_1 _3161_ (.A(_1421_),
    .X(_0158_));
 sky130_fd_sc_hd__or3_4 _3162_ (.A(_0720_),
    .B(_0727_),
    .C(_1409_),
    .X(_1422_));
 sky130_fd_sc_hd__or2_2 _3163_ (.A(_0921_),
    .B(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__mux2_1 _3164_ (.A0(_1381_),
    .A1(\tms1x00.RAM[108][0] ),
    .S(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_1 _3165_ (.A(_1424_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _3166_ (.A0(_1386_),
    .A1(\tms1x00.RAM[108][1] ),
    .S(_1423_),
    .X(_1425_));
 sky130_fd_sc_hd__clkbuf_1 _3167_ (.A(_1425_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _3168_ (.A0(_1388_),
    .A1(\tms1x00.RAM[108][2] ),
    .S(_1423_),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_1 _3169_ (.A(_1426_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _3170_ (.A0(_1390_),
    .A1(\tms1x00.RAM[108][3] ),
    .S(_1423_),
    .X(_1427_));
 sky130_fd_sc_hd__clkbuf_1 _3171_ (.A(_1427_),
    .X(_0162_));
 sky130_fd_sc_hd__or2_2 _3172_ (.A(_0921_),
    .B(_1288_),
    .X(_1428_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(_1381_),
    .A1(\tms1x00.RAM[107][0] ),
    .S(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__clkbuf_1 _3174_ (.A(_1429_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(_1386_),
    .A1(\tms1x00.RAM[107][1] ),
    .S(_1428_),
    .X(_1430_));
 sky130_fd_sc_hd__clkbuf_1 _3176_ (.A(_1430_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _3177_ (.A0(_1388_),
    .A1(\tms1x00.RAM[107][2] ),
    .S(_1428_),
    .X(_1431_));
 sky130_fd_sc_hd__clkbuf_1 _3178_ (.A(_1431_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _3179_ (.A0(_1390_),
    .A1(\tms1x00.RAM[107][3] ),
    .S(_1428_),
    .X(_1432_));
 sky130_fd_sc_hd__clkbuf_1 _3180_ (.A(_1432_),
    .X(_0166_));
 sky130_fd_sc_hd__or2_2 _3181_ (.A(_0921_),
    .B(_1416_),
    .X(_1433_));
 sky130_fd_sc_hd__mux2_1 _3182_ (.A0(_1381_),
    .A1(\tms1x00.RAM[106][0] ),
    .S(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_1 _3183_ (.A(_1434_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _3184_ (.A0(_1386_),
    .A1(\tms1x00.RAM[106][1] ),
    .S(_1433_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _3185_ (.A(_1435_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _3186_ (.A0(_1388_),
    .A1(\tms1x00.RAM[106][2] ),
    .S(_1433_),
    .X(_1436_));
 sky130_fd_sc_hd__clkbuf_1 _3187_ (.A(_1436_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _3188_ (.A0(_1390_),
    .A1(\tms1x00.RAM[106][3] ),
    .S(_1433_),
    .X(_1437_));
 sky130_fd_sc_hd__clkbuf_1 _3189_ (.A(_1437_),
    .X(_0170_));
 sky130_fd_sc_hd__or2_2 _3190_ (.A(_0921_),
    .B(_1255_),
    .X(_1438_));
 sky130_fd_sc_hd__mux2_1 _3191_ (.A0(_1381_),
    .A1(\tms1x00.RAM[105][0] ),
    .S(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__clkbuf_1 _3192_ (.A(_1439_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _3193_ (.A0(_1386_),
    .A1(\tms1x00.RAM[105][1] ),
    .S(_1438_),
    .X(_1440_));
 sky130_fd_sc_hd__clkbuf_1 _3194_ (.A(_1440_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _3195_ (.A0(_1388_),
    .A1(\tms1x00.RAM[105][2] ),
    .S(_1438_),
    .X(_1441_));
 sky130_fd_sc_hd__clkbuf_1 _3196_ (.A(_1441_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _3197_ (.A0(_1390_),
    .A1(\tms1x00.RAM[105][3] ),
    .S(_1438_),
    .X(_1442_));
 sky130_fd_sc_hd__clkbuf_1 _3198_ (.A(_1442_),
    .X(_0174_));
 sky130_fd_sc_hd__or2_2 _3199_ (.A(_1383_),
    .B(_1422_),
    .X(_1443_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(_1381_),
    .A1(\tms1x00.RAM[124][0] ),
    .S(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _3201_ (.A(_1444_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(_1386_),
    .A1(\tms1x00.RAM[124][1] ),
    .S(_1443_),
    .X(_1445_));
 sky130_fd_sc_hd__clkbuf_1 _3203_ (.A(_1445_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _3204_ (.A0(_1388_),
    .A1(\tms1x00.RAM[124][2] ),
    .S(_1443_),
    .X(_1446_));
 sky130_fd_sc_hd__clkbuf_1 _3205_ (.A(_1446_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _3206_ (.A0(_1390_),
    .A1(\tms1x00.RAM[124][3] ),
    .S(_1443_),
    .X(_1447_));
 sky130_fd_sc_hd__clkbuf_1 _3207_ (.A(_1447_),
    .X(_0178_));
 sky130_fd_sc_hd__nor2_4 _3208_ (.A(_1287_),
    .B(_1397_),
    .Y(_1448_));
 sky130_fd_sc_hd__mux2_1 _3209_ (.A0(\tms1x00.RAM[123][0] ),
    .A1(_1336_),
    .S(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__clkbuf_1 _3210_ (.A(_1449_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(\tms1x00.RAM[123][1] ),
    .A1(_1343_),
    .S(_1448_),
    .X(_1450_));
 sky130_fd_sc_hd__clkbuf_1 _3212_ (.A(_1450_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _3213_ (.A0(\tms1x00.RAM[123][2] ),
    .A1(_1346_),
    .S(_1448_),
    .X(_1451_));
 sky130_fd_sc_hd__clkbuf_1 _3214_ (.A(_1451_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(\tms1x00.RAM[123][3] ),
    .A1(_1349_),
    .S(_1448_),
    .X(_1452_));
 sky130_fd_sc_hd__clkbuf_1 _3216_ (.A(_1452_),
    .X(_0182_));
 sky130_fd_sc_hd__clkbuf_4 _3217_ (.A(_0919_),
    .X(_1453_));
 sky130_fd_sc_hd__or2_2 _3218_ (.A(_1383_),
    .B(_1416_),
    .X(_1454_));
 sky130_fd_sc_hd__mux2_1 _3219_ (.A0(_1453_),
    .A1(\tms1x00.RAM[122][0] ),
    .S(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_1 _3220_ (.A(_1455_),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_4 _3221_ (.A(_1031_),
    .X(_1456_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(_1456_),
    .A1(\tms1x00.RAM[122][1] ),
    .S(_1454_),
    .X(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _3223_ (.A(_1457_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_4 _3224_ (.A(_1132_),
    .X(_1458_));
 sky130_fd_sc_hd__mux2_1 _3225_ (.A0(_1458_),
    .A1(\tms1x00.RAM[122][2] ),
    .S(_1454_),
    .X(_1459_));
 sky130_fd_sc_hd__clkbuf_1 _3226_ (.A(_1459_),
    .X(_0185_));
 sky130_fd_sc_hd__clkbuf_4 _3227_ (.A(_1228_),
    .X(_1460_));
 sky130_fd_sc_hd__mux2_1 _3228_ (.A0(_1460_),
    .A1(\tms1x00.RAM[122][3] ),
    .S(_1454_),
    .X(_1461_));
 sky130_fd_sc_hd__clkbuf_1 _3229_ (.A(_1461_),
    .X(_0186_));
 sky130_fd_sc_hd__or2_2 _3230_ (.A(_1255_),
    .B(_1383_),
    .X(_1462_));
 sky130_fd_sc_hd__mux2_1 _3231_ (.A0(_1453_),
    .A1(\tms1x00.RAM[121][0] ),
    .S(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__clkbuf_1 _3232_ (.A(_1463_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _3233_ (.A0(_1456_),
    .A1(\tms1x00.RAM[121][1] ),
    .S(_1462_),
    .X(_1464_));
 sky130_fd_sc_hd__clkbuf_1 _3234_ (.A(_1464_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _3235_ (.A0(_1458_),
    .A1(\tms1x00.RAM[121][2] ),
    .S(_1462_),
    .X(_1465_));
 sky130_fd_sc_hd__clkbuf_1 _3236_ (.A(_1465_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _3237_ (.A0(_1460_),
    .A1(\tms1x00.RAM[121][3] ),
    .S(_1462_),
    .X(_1466_));
 sky130_fd_sc_hd__clkbuf_1 _3238_ (.A(_1466_),
    .X(_0190_));
 sky130_fd_sc_hd__or2_2 _3239_ (.A(_1309_),
    .B(_1383_),
    .X(_1467_));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(_1453_),
    .A1(\tms1x00.RAM[120][0] ),
    .S(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _3241_ (.A(_1468_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _3242_ (.A0(_1456_),
    .A1(\tms1x00.RAM[120][1] ),
    .S(_1467_),
    .X(_1469_));
 sky130_fd_sc_hd__clkbuf_1 _3243_ (.A(_1469_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _3244_ (.A0(_1458_),
    .A1(\tms1x00.RAM[120][2] ),
    .S(_1467_),
    .X(_1470_));
 sky130_fd_sc_hd__clkbuf_1 _3245_ (.A(_1470_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _3246_ (.A0(_1460_),
    .A1(\tms1x00.RAM[120][3] ),
    .S(_1467_),
    .X(_1471_));
 sky130_fd_sc_hd__clkbuf_1 _3247_ (.A(_1471_),
    .X(_0194_));
 sky130_fd_sc_hd__or2_1 _3248_ (.A(_0926_),
    .B(_1351_),
    .X(_1472_));
 sky130_fd_sc_hd__buf_2 _3249_ (.A(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__nor2_2 _3250_ (.A(_1287_),
    .B(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__mux2_1 _3251_ (.A0(\tms1x00.RAM[11][0] ),
    .A1(_1336_),
    .S(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__clkbuf_1 _3252_ (.A(_1475_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _3253_ (.A0(\tms1x00.RAM[11][1] ),
    .A1(_1343_),
    .S(_1474_),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_1 _3254_ (.A(_1476_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _3255_ (.A0(\tms1x00.RAM[11][2] ),
    .A1(_1346_),
    .S(_1474_),
    .X(_1477_));
 sky130_fd_sc_hd__clkbuf_1 _3256_ (.A(_1477_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _3257_ (.A0(\tms1x00.RAM[11][3] ),
    .A1(_1349_),
    .S(_1474_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_1 _3258_ (.A(_1478_),
    .X(_0198_));
 sky130_fd_sc_hd__nor2_2 _3259_ (.A(_1324_),
    .B(_1383_),
    .Y(_1479_));
 sky130_fd_sc_hd__mux2_1 _3260_ (.A0(\tms1x00.RAM[118][0] ),
    .A1(_1336_),
    .S(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__clkbuf_1 _3261_ (.A(_1480_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(\tms1x00.RAM[118][1] ),
    .A1(_1343_),
    .S(_1479_),
    .X(_1481_));
 sky130_fd_sc_hd__clkbuf_1 _3263_ (.A(_1481_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(\tms1x00.RAM[118][2] ),
    .A1(_1346_),
    .S(_1479_),
    .X(_1482_));
 sky130_fd_sc_hd__clkbuf_1 _3265_ (.A(_1482_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _3266_ (.A0(\tms1x00.RAM[118][3] ),
    .A1(_1349_),
    .S(_1479_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_1 _3267_ (.A(_1483_),
    .X(_0202_));
 sky130_fd_sc_hd__or2_2 _3268_ (.A(_1278_),
    .B(_1382_),
    .X(_1484_));
 sky130_fd_sc_hd__mux2_1 _3269_ (.A0(_1453_),
    .A1(\tms1x00.RAM[117][0] ),
    .S(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__clkbuf_1 _3270_ (.A(_1485_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _3271_ (.A0(_1456_),
    .A1(\tms1x00.RAM[117][1] ),
    .S(_1484_),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_1 _3272_ (.A(_1486_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _3273_ (.A0(_1458_),
    .A1(\tms1x00.RAM[117][2] ),
    .S(_1484_),
    .X(_1487_));
 sky130_fd_sc_hd__clkbuf_1 _3274_ (.A(_1487_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _3275_ (.A0(_1460_),
    .A1(\tms1x00.RAM[117][3] ),
    .S(_1484_),
    .X(_1488_));
 sky130_fd_sc_hd__clkbuf_1 _3276_ (.A(_1488_),
    .X(_0206_));
 sky130_fd_sc_hd__nor2_2 _3277_ (.A(_1339_),
    .B(_1383_),
    .Y(_1489_));
 sky130_fd_sc_hd__mux2_1 _3278_ (.A0(\tms1x00.RAM[116][0] ),
    .A1(_1336_),
    .S(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__clkbuf_1 _3279_ (.A(_1490_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _3280_ (.A0(\tms1x00.RAM[116][1] ),
    .A1(_1343_),
    .S(_1489_),
    .X(_1491_));
 sky130_fd_sc_hd__clkbuf_1 _3281_ (.A(_1491_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _3282_ (.A0(\tms1x00.RAM[116][2] ),
    .A1(_1346_),
    .S(_1489_),
    .X(_1492_));
 sky130_fd_sc_hd__clkbuf_1 _3283_ (.A(_1492_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _3284_ (.A0(\tms1x00.RAM[116][3] ),
    .A1(_1349_),
    .S(_1489_),
    .X(_1493_));
 sky130_fd_sc_hd__clkbuf_1 _3285_ (.A(_1493_),
    .X(_0210_));
 sky130_fd_sc_hd__or2_2 _3286_ (.A(_1233_),
    .B(_1382_),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_1 _3287_ (.A0(_1453_),
    .A1(\tms1x00.RAM[115][0] ),
    .S(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__clkbuf_1 _3288_ (.A(_1495_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _3289_ (.A0(_1456_),
    .A1(\tms1x00.RAM[115][1] ),
    .S(_1494_),
    .X(_1496_));
 sky130_fd_sc_hd__clkbuf_1 _3290_ (.A(_1496_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _3291_ (.A0(_1458_),
    .A1(\tms1x00.RAM[115][2] ),
    .S(_1494_),
    .X(_1497_));
 sky130_fd_sc_hd__clkbuf_1 _3292_ (.A(_1497_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _3293_ (.A0(_1460_),
    .A1(\tms1x00.RAM[115][3] ),
    .S(_1494_),
    .X(_1498_));
 sky130_fd_sc_hd__clkbuf_1 _3294_ (.A(_1498_),
    .X(_0214_));
 sky130_fd_sc_hd__or2_2 _3295_ (.A(_1383_),
    .B(_1410_),
    .X(_1499_));
 sky130_fd_sc_hd__mux2_1 _3296_ (.A0(_1453_),
    .A1(\tms1x00.RAM[126][0] ),
    .S(_1499_),
    .X(_1500_));
 sky130_fd_sc_hd__clkbuf_1 _3297_ (.A(_1500_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _3298_ (.A0(_1456_),
    .A1(\tms1x00.RAM[126][1] ),
    .S(_1499_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _3299_ (.A(_1501_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _3300_ (.A0(_1458_),
    .A1(\tms1x00.RAM[126][2] ),
    .S(_1499_),
    .X(_1502_));
 sky130_fd_sc_hd__clkbuf_1 _3301_ (.A(_1502_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _3302_ (.A0(_1460_),
    .A1(\tms1x00.RAM[126][3] ),
    .S(_1499_),
    .X(_1503_));
 sky130_fd_sc_hd__clkbuf_1 _3303_ (.A(_1503_),
    .X(_0218_));
 sky130_fd_sc_hd__nor2_2 _3304_ (.A(_0928_),
    .B(_1383_),
    .Y(_1504_));
 sky130_fd_sc_hd__mux2_1 _3305_ (.A0(\tms1x00.RAM[125][0] ),
    .A1(_1336_),
    .S(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__clkbuf_1 _3306_ (.A(_1505_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _3307_ (.A0(\tms1x00.RAM[125][1] ),
    .A1(_1343_),
    .S(_1504_),
    .X(_1506_));
 sky130_fd_sc_hd__clkbuf_1 _3308_ (.A(_1506_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _3309_ (.A0(\tms1x00.RAM[125][2] ),
    .A1(_1346_),
    .S(_1504_),
    .X(_1507_));
 sky130_fd_sc_hd__clkbuf_1 _3310_ (.A(_1507_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _3311_ (.A0(\tms1x00.RAM[125][3] ),
    .A1(_1349_),
    .S(_1504_),
    .X(_1508_));
 sky130_fd_sc_hd__clkbuf_1 _3312_ (.A(_1508_),
    .X(_0222_));
 sky130_fd_sc_hd__or2_2 _3313_ (.A(_1241_),
    .B(_1255_),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_1 _3314_ (.A0(_1453_),
    .A1(\tms1x00.RAM[25][0] ),
    .S(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_1 _3315_ (.A(_1510_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _3316_ (.A0(_1456_),
    .A1(\tms1x00.RAM[25][1] ),
    .S(_1509_),
    .X(_1511_));
 sky130_fd_sc_hd__clkbuf_1 _3317_ (.A(_1511_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _3318_ (.A0(_1458_),
    .A1(\tms1x00.RAM[25][2] ),
    .S(_1509_),
    .X(_1512_));
 sky130_fd_sc_hd__clkbuf_1 _3319_ (.A(_1512_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _3320_ (.A0(_1460_),
    .A1(\tms1x00.RAM[25][3] ),
    .S(_1509_),
    .X(_1513_));
 sky130_fd_sc_hd__clkbuf_1 _3321_ (.A(_1513_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_4 _3322_ (.A(_1335_),
    .X(_1514_));
 sky130_fd_sc_hd__nor2_2 _3323_ (.A(_1241_),
    .B(_1309_),
    .Y(_1515_));
 sky130_fd_sc_hd__mux2_1 _3324_ (.A0(\tms1x00.RAM[24][0] ),
    .A1(_1514_),
    .S(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__clkbuf_1 _3325_ (.A(_1516_),
    .X(_0227_));
 sky130_fd_sc_hd__clkbuf_4 _3326_ (.A(_1342_),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_1 _3327_ (.A0(\tms1x00.RAM[24][1] ),
    .A1(_1517_),
    .S(_1515_),
    .X(_1518_));
 sky130_fd_sc_hd__clkbuf_1 _3328_ (.A(_1518_),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_4 _3329_ (.A(_1345_),
    .X(_1519_));
 sky130_fd_sc_hd__mux2_1 _3330_ (.A0(\tms1x00.RAM[24][2] ),
    .A1(_1519_),
    .S(_1515_),
    .X(_1520_));
 sky130_fd_sc_hd__clkbuf_1 _3331_ (.A(_1520_),
    .X(_0229_));
 sky130_fd_sc_hd__clkbuf_4 _3332_ (.A(_1348_),
    .X(_1521_));
 sky130_fd_sc_hd__mux2_1 _3333_ (.A0(\tms1x00.RAM[24][3] ),
    .A1(_1521_),
    .S(_1515_),
    .X(_1522_));
 sky130_fd_sc_hd__clkbuf_1 _3334_ (.A(_1522_),
    .X(_0230_));
 sky130_fd_sc_hd__or2_2 _3335_ (.A(_1241_),
    .B(_1288_),
    .X(_1523_));
 sky130_fd_sc_hd__mux2_1 _3336_ (.A0(_1453_),
    .A1(\tms1x00.RAM[27][0] ),
    .S(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__clkbuf_1 _3337_ (.A(_1524_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _3338_ (.A0(_1456_),
    .A1(\tms1x00.RAM[27][1] ),
    .S(_1523_),
    .X(_1525_));
 sky130_fd_sc_hd__clkbuf_1 _3339_ (.A(_1525_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _3340_ (.A0(_1458_),
    .A1(\tms1x00.RAM[27][2] ),
    .S(_1523_),
    .X(_1526_));
 sky130_fd_sc_hd__clkbuf_1 _3341_ (.A(_1526_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _3342_ (.A0(_1460_),
    .A1(\tms1x00.RAM[27][3] ),
    .S(_1523_),
    .X(_1527_));
 sky130_fd_sc_hd__clkbuf_1 _3343_ (.A(_1527_),
    .X(_0234_));
 sky130_fd_sc_hd__or2_2 _3344_ (.A(_1241_),
    .B(_1416_),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _3345_ (.A0(_1453_),
    .A1(\tms1x00.RAM[26][0] ),
    .S(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__clkbuf_1 _3346_ (.A(_1529_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _3347_ (.A0(_1456_),
    .A1(\tms1x00.RAM[26][1] ),
    .S(_1528_),
    .X(_1530_));
 sky130_fd_sc_hd__clkbuf_1 _3348_ (.A(_1530_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _3349_ (.A0(_1458_),
    .A1(\tms1x00.RAM[26][2] ),
    .S(_1528_),
    .X(_1531_));
 sky130_fd_sc_hd__clkbuf_1 _3350_ (.A(_1531_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _3351_ (.A0(_1460_),
    .A1(\tms1x00.RAM[26][3] ),
    .S(_1528_),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_1 _3352_ (.A(_1532_),
    .X(_0238_));
 sky130_fd_sc_hd__or3b_4 _3353_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C_N(\tms1x00.ram_addr_buff[5] ),
    .X(_1533_));
 sky130_fd_sc_hd__buf_4 _3354_ (.A(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__nor2_2 _3355_ (.A(_1355_),
    .B(_1534_),
    .Y(_1535_));
 sky130_fd_sc_hd__mux2_1 _3356_ (.A0(\tms1x00.RAM[32][0] ),
    .A1(_1514_),
    .S(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__clkbuf_1 _3357_ (.A(_1536_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _3358_ (.A0(\tms1x00.RAM[32][1] ),
    .A1(_1517_),
    .S(_1535_),
    .X(_1537_));
 sky130_fd_sc_hd__clkbuf_1 _3359_ (.A(_1537_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _3360_ (.A0(\tms1x00.RAM[32][2] ),
    .A1(_1519_),
    .S(_1535_),
    .X(_1538_));
 sky130_fd_sc_hd__clkbuf_1 _3361_ (.A(_1538_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _3362_ (.A0(\tms1x00.RAM[32][3] ),
    .A1(_1521_),
    .S(_1535_),
    .X(_1539_));
 sky130_fd_sc_hd__clkbuf_1 _3363_ (.A(_1539_),
    .X(_0242_));
 sky130_fd_sc_hd__nor2_2 _3364_ (.A(_1241_),
    .B(_1403_),
    .Y(_1540_));
 sky130_fd_sc_hd__mux2_1 _3365_ (.A0(\tms1x00.RAM[31][0] ),
    .A1(_1514_),
    .S(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _3366_ (.A(_1541_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _3367_ (.A0(\tms1x00.RAM[31][1] ),
    .A1(_1517_),
    .S(_1540_),
    .X(_1542_));
 sky130_fd_sc_hd__clkbuf_1 _3368_ (.A(_1542_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _3369_ (.A0(\tms1x00.RAM[31][2] ),
    .A1(_1519_),
    .S(_1540_),
    .X(_1543_));
 sky130_fd_sc_hd__clkbuf_1 _3370_ (.A(_1543_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(\tms1x00.RAM[31][3] ),
    .A1(_1521_),
    .S(_1540_),
    .X(_1544_));
 sky130_fd_sc_hd__clkbuf_1 _3372_ (.A(_1544_),
    .X(_0246_));
 sky130_fd_sc_hd__or2_1 _3373_ (.A(_1240_),
    .B(_1410_),
    .X(_1545_));
 sky130_fd_sc_hd__mux2_1 _3374_ (.A0(_1453_),
    .A1(\tms1x00.RAM[30][0] ),
    .S(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__clkbuf_1 _3375_ (.A(_1546_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _3376_ (.A0(_1456_),
    .A1(\tms1x00.RAM[30][1] ),
    .S(_1545_),
    .X(_1547_));
 sky130_fd_sc_hd__clkbuf_1 _3377_ (.A(_1547_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _3378_ (.A0(_1458_),
    .A1(\tms1x00.RAM[30][2] ),
    .S(_1545_),
    .X(_1548_));
 sky130_fd_sc_hd__clkbuf_1 _3379_ (.A(_1548_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _3380_ (.A0(_1460_),
    .A1(\tms1x00.RAM[30][3] ),
    .S(_1545_),
    .X(_1549_));
 sky130_fd_sc_hd__clkbuf_1 _3381_ (.A(_1549_),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_4 _3382_ (.A(_0919_),
    .X(_1550_));
 sky130_fd_sc_hd__or2_2 _3383_ (.A(_1271_),
    .B(_1352_),
    .X(_1551_));
 sky130_fd_sc_hd__mux2_1 _3384_ (.A0(_1550_),
    .A1(\tms1x00.RAM[2][0] ),
    .S(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__clkbuf_1 _3385_ (.A(_1552_),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_4 _3386_ (.A(_1031_),
    .X(_1553_));
 sky130_fd_sc_hd__mux2_1 _3387_ (.A0(_1553_),
    .A1(\tms1x00.RAM[2][1] ),
    .S(_1551_),
    .X(_1554_));
 sky130_fd_sc_hd__clkbuf_1 _3388_ (.A(_1554_),
    .X(_0252_));
 sky130_fd_sc_hd__clkbuf_4 _3389_ (.A(_1132_),
    .X(_1555_));
 sky130_fd_sc_hd__mux2_1 _3390_ (.A0(_1555_),
    .A1(\tms1x00.RAM[2][2] ),
    .S(_1551_),
    .X(_1556_));
 sky130_fd_sc_hd__clkbuf_1 _3391_ (.A(_1556_),
    .X(_0253_));
 sky130_fd_sc_hd__clkbuf_4 _3392_ (.A(_1228_),
    .X(_1557_));
 sky130_fd_sc_hd__mux2_1 _3393_ (.A0(_1557_),
    .A1(\tms1x00.RAM[2][3] ),
    .S(_1551_),
    .X(_1558_));
 sky130_fd_sc_hd__clkbuf_1 _3394_ (.A(_1558_),
    .X(_0254_));
 sky130_fd_sc_hd__or2_2 _3395_ (.A(_1240_),
    .B(_1422_),
    .X(_1559_));
 sky130_fd_sc_hd__mux2_1 _3396_ (.A0(_1550_),
    .A1(\tms1x00.RAM[28][0] ),
    .S(_1559_),
    .X(_1560_));
 sky130_fd_sc_hd__clkbuf_1 _3397_ (.A(_1560_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _3398_ (.A0(_1553_),
    .A1(\tms1x00.RAM[28][1] ),
    .S(_1559_),
    .X(_1561_));
 sky130_fd_sc_hd__clkbuf_1 _3399_ (.A(_1561_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _3400_ (.A0(_1555_),
    .A1(\tms1x00.RAM[28][2] ),
    .S(_1559_),
    .X(_1562_));
 sky130_fd_sc_hd__clkbuf_1 _3401_ (.A(_1562_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _3402_ (.A0(_1557_),
    .A1(\tms1x00.RAM[28][3] ),
    .S(_1559_),
    .X(_1563_));
 sky130_fd_sc_hd__clkbuf_1 _3403_ (.A(_1563_),
    .X(_0258_));
 sky130_fd_sc_hd__nor2_2 _3404_ (.A(_1339_),
    .B(_1534_),
    .Y(_1564_));
 sky130_fd_sc_hd__mux2_1 _3405_ (.A0(\tms1x00.RAM[36][0] ),
    .A1(_1514_),
    .S(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__clkbuf_1 _3406_ (.A(_1565_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _3407_ (.A0(\tms1x00.RAM[36][1] ),
    .A1(_1517_),
    .S(_1564_),
    .X(_1566_));
 sky130_fd_sc_hd__clkbuf_1 _3408_ (.A(_1566_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _3409_ (.A0(\tms1x00.RAM[36][2] ),
    .A1(_1519_),
    .S(_1564_),
    .X(_1567_));
 sky130_fd_sc_hd__clkbuf_1 _3410_ (.A(_1567_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _3411_ (.A0(\tms1x00.RAM[36][3] ),
    .A1(_1521_),
    .S(_1564_),
    .X(_1568_));
 sky130_fd_sc_hd__clkbuf_1 _3412_ (.A(_1568_),
    .X(_0262_));
 sky130_fd_sc_hd__nor2_2 _3413_ (.A(_1233_),
    .B(_1534_),
    .Y(_1569_));
 sky130_fd_sc_hd__mux2_1 _3414_ (.A0(\tms1x00.RAM[35][0] ),
    .A1(_1514_),
    .S(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__clkbuf_1 _3415_ (.A(_1570_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _3416_ (.A0(\tms1x00.RAM[35][1] ),
    .A1(_1517_),
    .S(_1569_),
    .X(_1571_));
 sky130_fd_sc_hd__clkbuf_1 _3417_ (.A(_1571_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _3418_ (.A0(\tms1x00.RAM[35][2] ),
    .A1(_1519_),
    .S(_1569_),
    .X(_1572_));
 sky130_fd_sc_hd__clkbuf_1 _3419_ (.A(_1572_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _3420_ (.A0(\tms1x00.RAM[35][3] ),
    .A1(_1521_),
    .S(_1569_),
    .X(_1573_));
 sky130_fd_sc_hd__clkbuf_1 _3421_ (.A(_1573_),
    .X(_0266_));
 sky130_fd_sc_hd__or2_2 _3422_ (.A(_1271_),
    .B(_1534_),
    .X(_1574_));
 sky130_fd_sc_hd__mux2_1 _3423_ (.A0(_1550_),
    .A1(\tms1x00.RAM[34][0] ),
    .S(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__clkbuf_1 _3424_ (.A(_1575_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _3425_ (.A0(_1553_),
    .A1(\tms1x00.RAM[34][1] ),
    .S(_1574_),
    .X(_1576_));
 sky130_fd_sc_hd__clkbuf_1 _3426_ (.A(_1576_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _3427_ (.A0(_1555_),
    .A1(\tms1x00.RAM[34][2] ),
    .S(_1574_),
    .X(_1577_));
 sky130_fd_sc_hd__clkbuf_1 _3428_ (.A(_1577_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _3429_ (.A0(_1557_),
    .A1(\tms1x00.RAM[34][3] ),
    .S(_1574_),
    .X(_1578_));
 sky130_fd_sc_hd__clkbuf_1 _3430_ (.A(_1578_),
    .X(_0270_));
 sky130_fd_sc_hd__or2_2 _3431_ (.A(_1243_),
    .B(_1533_),
    .X(_1579_));
 sky130_fd_sc_hd__mux2_1 _3432_ (.A0(_1550_),
    .A1(\tms1x00.RAM[33][0] ),
    .S(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__clkbuf_1 _3433_ (.A(_1580_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _3434_ (.A0(_1553_),
    .A1(\tms1x00.RAM[33][1] ),
    .S(_1579_),
    .X(_1581_));
 sky130_fd_sc_hd__clkbuf_1 _3435_ (.A(_1581_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _3436_ (.A0(_1555_),
    .A1(\tms1x00.RAM[33][2] ),
    .S(_1579_),
    .X(_1582_));
 sky130_fd_sc_hd__clkbuf_1 _3437_ (.A(_1582_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(_1557_),
    .A1(\tms1x00.RAM[33][3] ),
    .S(_1579_),
    .X(_1583_));
 sky130_fd_sc_hd__clkbuf_1 _3439_ (.A(_1583_),
    .X(_0274_));
 sky130_fd_sc_hd__or2_2 _3440_ (.A(_1255_),
    .B(_1533_),
    .X(_1584_));
 sky130_fd_sc_hd__mux2_1 _3441_ (.A0(_1550_),
    .A1(\tms1x00.RAM[41][0] ),
    .S(_1584_),
    .X(_1585_));
 sky130_fd_sc_hd__clkbuf_1 _3442_ (.A(_1585_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _3443_ (.A0(_1553_),
    .A1(\tms1x00.RAM[41][1] ),
    .S(_1584_),
    .X(_1586_));
 sky130_fd_sc_hd__clkbuf_1 _3444_ (.A(_1586_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _3445_ (.A0(_1555_),
    .A1(\tms1x00.RAM[41][2] ),
    .S(_1584_),
    .X(_1587_));
 sky130_fd_sc_hd__clkbuf_1 _3446_ (.A(_1587_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _3447_ (.A0(_1557_),
    .A1(\tms1x00.RAM[41][3] ),
    .S(_1584_),
    .X(_1588_));
 sky130_fd_sc_hd__clkbuf_1 _3448_ (.A(_1588_),
    .X(_0278_));
 sky130_fd_sc_hd__nor2_2 _3449_ (.A(_1309_),
    .B(_1534_),
    .Y(_1589_));
 sky130_fd_sc_hd__mux2_1 _3450_ (.A0(\tms1x00.RAM[40][0] ),
    .A1(_1514_),
    .S(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__clkbuf_1 _3451_ (.A(_1590_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _3452_ (.A0(\tms1x00.RAM[40][1] ),
    .A1(_1517_),
    .S(_1589_),
    .X(_1591_));
 sky130_fd_sc_hd__clkbuf_1 _3453_ (.A(_1591_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _3454_ (.A0(\tms1x00.RAM[40][2] ),
    .A1(_1519_),
    .S(_1589_),
    .X(_1592_));
 sky130_fd_sc_hd__clkbuf_1 _3455_ (.A(_1592_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _3456_ (.A0(\tms1x00.RAM[40][3] ),
    .A1(_1521_),
    .S(_1589_),
    .X(_1593_));
 sky130_fd_sc_hd__clkbuf_1 _3457_ (.A(_1593_),
    .X(_0282_));
 sky130_fd_sc_hd__nor2_2 _3458_ (.A(_1233_),
    .B(_1352_),
    .Y(_1594_));
 sky130_fd_sc_hd__mux2_1 _3459_ (.A0(\tms1x00.RAM[3][0] ),
    .A1(_1514_),
    .S(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _3460_ (.A(_1595_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _3461_ (.A0(\tms1x00.RAM[3][1] ),
    .A1(_1517_),
    .S(_1594_),
    .X(_1596_));
 sky130_fd_sc_hd__clkbuf_1 _3462_ (.A(_1596_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _3463_ (.A0(\tms1x00.RAM[3][2] ),
    .A1(_1519_),
    .S(_1594_),
    .X(_1597_));
 sky130_fd_sc_hd__clkbuf_1 _3464_ (.A(_1597_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _3465_ (.A0(\tms1x00.RAM[3][3] ),
    .A1(_1521_),
    .S(_1594_),
    .X(_1598_));
 sky130_fd_sc_hd__clkbuf_1 _3466_ (.A(_1598_),
    .X(_0286_));
 sky130_fd_sc_hd__nor2_2 _3467_ (.A(_1324_),
    .B(_1534_),
    .Y(_1599_));
 sky130_fd_sc_hd__mux2_1 _3468_ (.A0(\tms1x00.RAM[38][0] ),
    .A1(_1514_),
    .S(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__clkbuf_1 _3469_ (.A(_1600_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _3470_ (.A0(\tms1x00.RAM[38][1] ),
    .A1(_1517_),
    .S(_1599_),
    .X(_1601_));
 sky130_fd_sc_hd__clkbuf_1 _3471_ (.A(_1601_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _3472_ (.A0(\tms1x00.RAM[38][2] ),
    .A1(_1519_),
    .S(_1599_),
    .X(_1602_));
 sky130_fd_sc_hd__clkbuf_1 _3473_ (.A(_1602_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _3474_ (.A0(\tms1x00.RAM[38][3] ),
    .A1(_1521_),
    .S(_1599_),
    .X(_1603_));
 sky130_fd_sc_hd__clkbuf_1 _3475_ (.A(_1603_),
    .X(_0290_));
 sky130_fd_sc_hd__or2_2 _3476_ (.A(_1278_),
    .B(_1533_),
    .X(_1604_));
 sky130_fd_sc_hd__mux2_1 _3477_ (.A0(_1550_),
    .A1(\tms1x00.RAM[37][0] ),
    .S(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__clkbuf_1 _3478_ (.A(_1605_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _3479_ (.A0(_1553_),
    .A1(\tms1x00.RAM[37][1] ),
    .S(_1604_),
    .X(_1606_));
 sky130_fd_sc_hd__clkbuf_1 _3480_ (.A(_1606_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _3481_ (.A0(_1555_),
    .A1(\tms1x00.RAM[37][2] ),
    .S(_1604_),
    .X(_1607_));
 sky130_fd_sc_hd__clkbuf_1 _3482_ (.A(_1607_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _3483_ (.A0(_1557_),
    .A1(\tms1x00.RAM[37][3] ),
    .S(_1604_),
    .X(_1608_));
 sky130_fd_sc_hd__clkbuf_1 _3484_ (.A(_1608_),
    .X(_0294_));
 sky130_fd_sc_hd__nor2_2 _3485_ (.A(_0928_),
    .B(_1534_),
    .Y(_1609_));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(\tms1x00.RAM[45][0] ),
    .A1(_1514_),
    .S(_1609_),
    .X(_1610_));
 sky130_fd_sc_hd__clkbuf_1 _3487_ (.A(_1610_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _3488_ (.A0(\tms1x00.RAM[45][1] ),
    .A1(_1517_),
    .S(_1609_),
    .X(_1611_));
 sky130_fd_sc_hd__clkbuf_1 _3489_ (.A(_1611_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _3490_ (.A0(\tms1x00.RAM[45][2] ),
    .A1(_1519_),
    .S(_1609_),
    .X(_1612_));
 sky130_fd_sc_hd__clkbuf_1 _3491_ (.A(_1612_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _3492_ (.A0(\tms1x00.RAM[45][3] ),
    .A1(_1521_),
    .S(_1609_),
    .X(_1613_));
 sky130_fd_sc_hd__clkbuf_1 _3493_ (.A(_1613_),
    .X(_0298_));
 sky130_fd_sc_hd__or2_2 _3494_ (.A(_1422_),
    .B(_1533_),
    .X(_1614_));
 sky130_fd_sc_hd__mux2_1 _3495_ (.A0(_1550_),
    .A1(\tms1x00.RAM[44][0] ),
    .S(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__clkbuf_1 _3496_ (.A(_1615_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _3497_ (.A0(_1553_),
    .A1(\tms1x00.RAM[44][1] ),
    .S(_1614_),
    .X(_1616_));
 sky130_fd_sc_hd__clkbuf_1 _3498_ (.A(_1616_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _3499_ (.A0(_1555_),
    .A1(\tms1x00.RAM[44][2] ),
    .S(_1614_),
    .X(_1617_));
 sky130_fd_sc_hd__clkbuf_1 _3500_ (.A(_1617_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _3501_ (.A0(_1557_),
    .A1(\tms1x00.RAM[44][3] ),
    .S(_1614_),
    .X(_1618_));
 sky130_fd_sc_hd__clkbuf_1 _3502_ (.A(_1618_),
    .X(_0302_));
 sky130_fd_sc_hd__nor2_2 _3503_ (.A(_1288_),
    .B(_1534_),
    .Y(_1619_));
 sky130_fd_sc_hd__mux2_1 _3504_ (.A0(\tms1x00.RAM[43][0] ),
    .A1(_1514_),
    .S(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__clkbuf_1 _3505_ (.A(_1620_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _3506_ (.A0(\tms1x00.RAM[43][1] ),
    .A1(_1517_),
    .S(_1619_),
    .X(_1621_));
 sky130_fd_sc_hd__clkbuf_1 _3507_ (.A(_1621_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _3508_ (.A0(\tms1x00.RAM[43][2] ),
    .A1(_1519_),
    .S(_1619_),
    .X(_1622_));
 sky130_fd_sc_hd__clkbuf_1 _3509_ (.A(_1622_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _3510_ (.A0(\tms1x00.RAM[43][3] ),
    .A1(_1521_),
    .S(_1619_),
    .X(_1623_));
 sky130_fd_sc_hd__clkbuf_1 _3511_ (.A(_1623_),
    .X(_0306_));
 sky130_fd_sc_hd__or2_2 _3512_ (.A(_1416_),
    .B(_1533_),
    .X(_1624_));
 sky130_fd_sc_hd__mux2_1 _3513_ (.A0(_1550_),
    .A1(\tms1x00.RAM[42][0] ),
    .S(_1624_),
    .X(_1625_));
 sky130_fd_sc_hd__clkbuf_1 _3514_ (.A(_1625_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(_1553_),
    .A1(\tms1x00.RAM[42][1] ),
    .S(_1624_),
    .X(_1626_));
 sky130_fd_sc_hd__clkbuf_1 _3516_ (.A(_1626_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _3517_ (.A0(_1555_),
    .A1(\tms1x00.RAM[42][2] ),
    .S(_1624_),
    .X(_1627_));
 sky130_fd_sc_hd__clkbuf_1 _3518_ (.A(_1627_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _3519_ (.A0(_1557_),
    .A1(\tms1x00.RAM[42][3] ),
    .S(_1624_),
    .X(_1628_));
 sky130_fd_sc_hd__clkbuf_1 _3520_ (.A(_1628_),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_4 _3521_ (.A(_0919_),
    .X(_1629_));
 sky130_fd_sc_hd__nor2_2 _3522_ (.A(_1337_),
    .B(_1473_),
    .Y(_1630_));
 sky130_fd_sc_hd__mux2_1 _3523_ (.A0(\tms1x00.RAM[4][0] ),
    .A1(_1629_),
    .S(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__clkbuf_1 _3524_ (.A(_1631_),
    .X(_0311_));
 sky130_fd_sc_hd__clkbuf_4 _3525_ (.A(_1031_),
    .X(_1632_));
 sky130_fd_sc_hd__mux2_1 _3526_ (.A0(\tms1x00.RAM[4][1] ),
    .A1(_1632_),
    .S(_1630_),
    .X(_1633_));
 sky130_fd_sc_hd__clkbuf_1 _3527_ (.A(_1633_),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_4 _3528_ (.A(_1132_),
    .X(_1634_));
 sky130_fd_sc_hd__mux2_1 _3529_ (.A0(\tms1x00.RAM[4][2] ),
    .A1(_1634_),
    .S(_1630_),
    .X(_1635_));
 sky130_fd_sc_hd__clkbuf_1 _3530_ (.A(_1635_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_4 _3531_ (.A(_1228_),
    .X(_1636_));
 sky130_fd_sc_hd__mux2_1 _3532_ (.A0(\tms1x00.RAM[4][3] ),
    .A1(_1636_),
    .S(_1630_),
    .X(_1637_));
 sky130_fd_sc_hd__clkbuf_1 _3533_ (.A(_1637_),
    .X(_0314_));
 sky130_fd_sc_hd__nor2_2 _3534_ (.A(_1285_),
    .B(_1355_),
    .Y(_1638_));
 sky130_fd_sc_hd__mux2_1 _3535_ (.A0(\tms1x00.RAM[48][0] ),
    .A1(_1629_),
    .S(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__clkbuf_1 _3536_ (.A(_1639_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _3537_ (.A0(\tms1x00.RAM[48][1] ),
    .A1(_1632_),
    .S(_1638_),
    .X(_1640_));
 sky130_fd_sc_hd__clkbuf_1 _3538_ (.A(_1640_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _3539_ (.A0(\tms1x00.RAM[48][2] ),
    .A1(_1634_),
    .S(_1638_),
    .X(_1641_));
 sky130_fd_sc_hd__clkbuf_1 _3540_ (.A(_1641_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _3541_ (.A0(\tms1x00.RAM[48][3] ),
    .A1(_1636_),
    .S(_1638_),
    .X(_1642_));
 sky130_fd_sc_hd__clkbuf_1 _3542_ (.A(_1642_),
    .X(_0318_));
 sky130_fd_sc_hd__nor2_2 _3543_ (.A(_1403_),
    .B(_1534_),
    .Y(_1643_));
 sky130_fd_sc_hd__mux2_1 _3544_ (.A0(\tms1x00.RAM[47][0] ),
    .A1(_1629_),
    .S(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__clkbuf_1 _3545_ (.A(_1644_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _3546_ (.A0(\tms1x00.RAM[47][1] ),
    .A1(_1632_),
    .S(_1643_),
    .X(_1645_));
 sky130_fd_sc_hd__clkbuf_1 _3547_ (.A(_1645_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _3548_ (.A0(\tms1x00.RAM[47][2] ),
    .A1(_1634_),
    .S(_1643_),
    .X(_1646_));
 sky130_fd_sc_hd__clkbuf_1 _3549_ (.A(_1646_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _3550_ (.A0(\tms1x00.RAM[47][3] ),
    .A1(_1636_),
    .S(_1643_),
    .X(_1647_));
 sky130_fd_sc_hd__clkbuf_1 _3551_ (.A(_1647_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_2 _3552_ (.A(_1410_),
    .B(_1533_),
    .X(_1648_));
 sky130_fd_sc_hd__mux2_1 _3553_ (.A0(_1550_),
    .A1(\tms1x00.RAM[46][0] ),
    .S(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__clkbuf_1 _3554_ (.A(_1649_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _3555_ (.A0(_1553_),
    .A1(\tms1x00.RAM[46][1] ),
    .S(_1648_),
    .X(_1650_));
 sky130_fd_sc_hd__clkbuf_1 _3556_ (.A(_1650_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _3557_ (.A0(_1555_),
    .A1(\tms1x00.RAM[46][2] ),
    .S(_1648_),
    .X(_1651_));
 sky130_fd_sc_hd__clkbuf_1 _3558_ (.A(_1651_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _3559_ (.A0(_1557_),
    .A1(\tms1x00.RAM[46][3] ),
    .S(_1648_),
    .X(_1652_));
 sky130_fd_sc_hd__clkbuf_1 _3560_ (.A(_1652_),
    .X(_0326_));
 sky130_fd_sc_hd__nor2_2 _3561_ (.A(_1285_),
    .B(_1324_),
    .Y(_1653_));
 sky130_fd_sc_hd__mux2_1 _3562_ (.A0(\tms1x00.RAM[54][0] ),
    .A1(_1629_),
    .S(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__clkbuf_1 _3563_ (.A(_1654_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _3564_ (.A0(\tms1x00.RAM[54][1] ),
    .A1(_1632_),
    .S(_1653_),
    .X(_1655_));
 sky130_fd_sc_hd__clkbuf_1 _3565_ (.A(_1655_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _3566_ (.A0(\tms1x00.RAM[54][2] ),
    .A1(_1634_),
    .S(_1653_),
    .X(_1656_));
 sky130_fd_sc_hd__clkbuf_1 _3567_ (.A(_1656_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _3568_ (.A0(\tms1x00.RAM[54][3] ),
    .A1(_1636_),
    .S(_1653_),
    .X(_1657_));
 sky130_fd_sc_hd__clkbuf_1 _3569_ (.A(_1657_),
    .X(_0330_));
 sky130_fd_sc_hd__or2_2 _3570_ (.A(_1278_),
    .B(_1284_),
    .X(_1658_));
 sky130_fd_sc_hd__mux2_1 _3571_ (.A0(_1550_),
    .A1(\tms1x00.RAM[53][0] ),
    .S(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__clkbuf_1 _3572_ (.A(_1659_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _3573_ (.A0(_1553_),
    .A1(\tms1x00.RAM[53][1] ),
    .S(_1658_),
    .X(_1660_));
 sky130_fd_sc_hd__clkbuf_1 _3574_ (.A(_1660_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _3575_ (.A0(_1555_),
    .A1(\tms1x00.RAM[53][2] ),
    .S(_1658_),
    .X(_1661_));
 sky130_fd_sc_hd__clkbuf_1 _3576_ (.A(_1661_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _3577_ (.A0(_1557_),
    .A1(\tms1x00.RAM[53][3] ),
    .S(_1658_),
    .X(_1662_));
 sky130_fd_sc_hd__clkbuf_1 _3578_ (.A(_1662_),
    .X(_0334_));
 sky130_fd_sc_hd__nor2_2 _3579_ (.A(_1285_),
    .B(_1339_),
    .Y(_1663_));
 sky130_fd_sc_hd__mux2_1 _3580_ (.A0(\tms1x00.RAM[52][0] ),
    .A1(_1629_),
    .S(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__clkbuf_1 _3581_ (.A(_1664_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _3582_ (.A0(\tms1x00.RAM[52][1] ),
    .A1(_1632_),
    .S(_1663_),
    .X(_1665_));
 sky130_fd_sc_hd__clkbuf_1 _3583_ (.A(_1665_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _3584_ (.A0(\tms1x00.RAM[52][2] ),
    .A1(_1634_),
    .S(_1663_),
    .X(_1666_));
 sky130_fd_sc_hd__clkbuf_1 _3585_ (.A(_1666_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _3586_ (.A0(\tms1x00.RAM[52][3] ),
    .A1(_1636_),
    .S(_1663_),
    .X(_1667_));
 sky130_fd_sc_hd__clkbuf_1 _3587_ (.A(_1667_),
    .X(_0338_));
 sky130_fd_sc_hd__nor2_2 _3588_ (.A(_1233_),
    .B(_1285_),
    .Y(_1668_));
 sky130_fd_sc_hd__mux2_1 _3589_ (.A0(\tms1x00.RAM[51][0] ),
    .A1(_1629_),
    .S(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__clkbuf_1 _3590_ (.A(_1669_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _3591_ (.A0(\tms1x00.RAM[51][1] ),
    .A1(_1632_),
    .S(_1668_),
    .X(_1670_));
 sky130_fd_sc_hd__clkbuf_1 _3592_ (.A(_1670_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _3593_ (.A0(\tms1x00.RAM[51][2] ),
    .A1(_1634_),
    .S(_1668_),
    .X(_1671_));
 sky130_fd_sc_hd__clkbuf_1 _3594_ (.A(_1671_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _3595_ (.A0(\tms1x00.RAM[51][3] ),
    .A1(_1636_),
    .S(_1668_),
    .X(_1672_));
 sky130_fd_sc_hd__clkbuf_1 _3596_ (.A(_1672_),
    .X(_0342_));
 sky130_fd_sc_hd__buf_2 _3597_ (.A(_0919_),
    .X(_1673_));
 sky130_fd_sc_hd__or2_2 _3598_ (.A(_1271_),
    .B(_1284_),
    .X(_1674_));
 sky130_fd_sc_hd__mux2_1 _3599_ (.A0(_1673_),
    .A1(\tms1x00.RAM[50][0] ),
    .S(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__clkbuf_1 _3600_ (.A(_1675_),
    .X(_0343_));
 sky130_fd_sc_hd__buf_2 _3601_ (.A(_1031_),
    .X(_1676_));
 sky130_fd_sc_hd__mux2_1 _3602_ (.A0(_1676_),
    .A1(\tms1x00.RAM[50][1] ),
    .S(_1674_),
    .X(_1677_));
 sky130_fd_sc_hd__clkbuf_1 _3603_ (.A(_1677_),
    .X(_0344_));
 sky130_fd_sc_hd__buf_2 _3604_ (.A(_1132_),
    .X(_1678_));
 sky130_fd_sc_hd__mux2_1 _3605_ (.A0(_1678_),
    .A1(\tms1x00.RAM[50][2] ),
    .S(_1674_),
    .X(_1679_));
 sky130_fd_sc_hd__clkbuf_1 _3606_ (.A(_1679_),
    .X(_0345_));
 sky130_fd_sc_hd__buf_2 _3607_ (.A(_1228_),
    .X(_1680_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(_1680_),
    .A1(\tms1x00.RAM[50][3] ),
    .S(_1674_),
    .X(_1681_));
 sky130_fd_sc_hd__clkbuf_1 _3609_ (.A(_1681_),
    .X(_0346_));
 sky130_fd_sc_hd__or2_2 _3610_ (.A(_1285_),
    .B(_1416_),
    .X(_1682_));
 sky130_fd_sc_hd__mux2_1 _3611_ (.A0(_1673_),
    .A1(\tms1x00.RAM[58][0] ),
    .S(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__clkbuf_1 _3612_ (.A(_1683_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _3613_ (.A0(_1676_),
    .A1(\tms1x00.RAM[58][1] ),
    .S(_1682_),
    .X(_1684_));
 sky130_fd_sc_hd__clkbuf_1 _3614_ (.A(_1684_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _3615_ (.A0(_1678_),
    .A1(\tms1x00.RAM[58][2] ),
    .S(_1682_),
    .X(_1685_));
 sky130_fd_sc_hd__clkbuf_1 _3616_ (.A(_1685_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _3617_ (.A0(_1680_),
    .A1(\tms1x00.RAM[58][3] ),
    .S(_1682_),
    .X(_1686_));
 sky130_fd_sc_hd__clkbuf_1 _3618_ (.A(_1686_),
    .X(_0350_));
 sky130_fd_sc_hd__or2_2 _3619_ (.A(_1255_),
    .B(_1284_),
    .X(_1687_));
 sky130_fd_sc_hd__mux2_1 _3620_ (.A0(_1673_),
    .A1(\tms1x00.RAM[57][0] ),
    .S(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__clkbuf_1 _3621_ (.A(_1688_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _3622_ (.A0(_1676_),
    .A1(\tms1x00.RAM[57][1] ),
    .S(_1687_),
    .X(_1689_));
 sky130_fd_sc_hd__clkbuf_1 _3623_ (.A(_1689_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _3624_ (.A0(_1678_),
    .A1(\tms1x00.RAM[57][2] ),
    .S(_1687_),
    .X(_1690_));
 sky130_fd_sc_hd__clkbuf_1 _3625_ (.A(_1690_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _3626_ (.A0(_1680_),
    .A1(\tms1x00.RAM[57][3] ),
    .S(_1687_),
    .X(_1691_));
 sky130_fd_sc_hd__clkbuf_1 _3627_ (.A(_1691_),
    .X(_0354_));
 sky130_fd_sc_hd__nor2_2 _3628_ (.A(_1285_),
    .B(_1309_),
    .Y(_1692_));
 sky130_fd_sc_hd__mux2_1 _3629_ (.A0(\tms1x00.RAM[56][0] ),
    .A1(_1629_),
    .S(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__clkbuf_1 _3630_ (.A(_1693_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _3631_ (.A0(\tms1x00.RAM[56][1] ),
    .A1(_1632_),
    .S(_1692_),
    .X(_1694_));
 sky130_fd_sc_hd__clkbuf_1 _3632_ (.A(_1694_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _3633_ (.A0(\tms1x00.RAM[56][2] ),
    .A1(_1634_),
    .S(_1692_),
    .X(_1695_));
 sky130_fd_sc_hd__clkbuf_1 _3634_ (.A(_1695_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _3635_ (.A0(\tms1x00.RAM[56][3] ),
    .A1(_1636_),
    .S(_1692_),
    .X(_1696_));
 sky130_fd_sc_hd__clkbuf_1 _3636_ (.A(_1696_),
    .X(_0358_));
 sky130_fd_sc_hd__or2_2 _3637_ (.A(_1242_),
    .B(_1316_),
    .X(_1697_));
 sky130_fd_sc_hd__nor2_2 _3638_ (.A(_1285_),
    .B(_1697_),
    .Y(_1698_));
 sky130_fd_sc_hd__mux2_1 _3639_ (.A0(\tms1x00.RAM[55][0] ),
    .A1(_1629_),
    .S(_1698_),
    .X(_1699_));
 sky130_fd_sc_hd__clkbuf_1 _3640_ (.A(_1699_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _3641_ (.A0(\tms1x00.RAM[55][1] ),
    .A1(_1632_),
    .S(_1698_),
    .X(_1700_));
 sky130_fd_sc_hd__clkbuf_1 _3642_ (.A(_1700_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _3643_ (.A0(\tms1x00.RAM[55][2] ),
    .A1(_1634_),
    .S(_1698_),
    .X(_1701_));
 sky130_fd_sc_hd__clkbuf_1 _3644_ (.A(_1701_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _3645_ (.A0(\tms1x00.RAM[55][3] ),
    .A1(_1636_),
    .S(_1698_),
    .X(_1702_));
 sky130_fd_sc_hd__clkbuf_1 _3646_ (.A(_1702_),
    .X(_0362_));
 sky130_fd_sc_hd__or2_2 _3647_ (.A(_1285_),
    .B(_1410_),
    .X(_1703_));
 sky130_fd_sc_hd__mux2_1 _3648_ (.A0(_1673_),
    .A1(\tms1x00.RAM[62][0] ),
    .S(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__clkbuf_1 _3649_ (.A(_1704_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _3650_ (.A0(_1676_),
    .A1(\tms1x00.RAM[62][1] ),
    .S(_1703_),
    .X(_1705_));
 sky130_fd_sc_hd__clkbuf_1 _3651_ (.A(_1705_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _3652_ (.A0(_1678_),
    .A1(\tms1x00.RAM[62][2] ),
    .S(_1703_),
    .X(_1706_));
 sky130_fd_sc_hd__clkbuf_1 _3653_ (.A(_1706_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _3654_ (.A0(_1680_),
    .A1(\tms1x00.RAM[62][3] ),
    .S(_1703_),
    .X(_1707_));
 sky130_fd_sc_hd__clkbuf_1 _3655_ (.A(_1707_),
    .X(_0366_));
 sky130_fd_sc_hd__nor2_2 _3656_ (.A(_0928_),
    .B(_1285_),
    .Y(_1708_));
 sky130_fd_sc_hd__mux2_1 _3657_ (.A0(\tms1x00.RAM[61][0] ),
    .A1(_1629_),
    .S(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__clkbuf_1 _3658_ (.A(_1709_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _3659_ (.A0(\tms1x00.RAM[61][1] ),
    .A1(_1632_),
    .S(_1708_),
    .X(_1710_));
 sky130_fd_sc_hd__clkbuf_1 _3660_ (.A(_1710_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _3661_ (.A0(\tms1x00.RAM[61][2] ),
    .A1(_1634_),
    .S(_1708_),
    .X(_1711_));
 sky130_fd_sc_hd__clkbuf_1 _3662_ (.A(_1711_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _3663_ (.A0(\tms1x00.RAM[61][3] ),
    .A1(_1636_),
    .S(_1708_),
    .X(_1712_));
 sky130_fd_sc_hd__clkbuf_1 _3664_ (.A(_1712_),
    .X(_0370_));
 sky130_fd_sc_hd__or2_2 _3665_ (.A(_1284_),
    .B(_1422_),
    .X(_1713_));
 sky130_fd_sc_hd__mux2_1 _3666_ (.A0(_1673_),
    .A1(\tms1x00.RAM[60][0] ),
    .S(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__clkbuf_1 _3667_ (.A(_1714_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _3668_ (.A0(_1676_),
    .A1(\tms1x00.RAM[60][1] ),
    .S(_1713_),
    .X(_1715_));
 sky130_fd_sc_hd__clkbuf_1 _3669_ (.A(_1715_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _3670_ (.A0(_1678_),
    .A1(\tms1x00.RAM[60][2] ),
    .S(_1713_),
    .X(_1716_));
 sky130_fd_sc_hd__clkbuf_1 _3671_ (.A(_1716_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _3672_ (.A0(_1680_),
    .A1(\tms1x00.RAM[60][3] ),
    .S(_1713_),
    .X(_1717_));
 sky130_fd_sc_hd__clkbuf_1 _3673_ (.A(_1717_),
    .X(_0374_));
 sky130_fd_sc_hd__or2_2 _3674_ (.A(_1278_),
    .B(_1352_),
    .X(_1718_));
 sky130_fd_sc_hd__mux2_1 _3675_ (.A0(_1673_),
    .A1(\tms1x00.RAM[5][0] ),
    .S(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__clkbuf_1 _3676_ (.A(_1719_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _3677_ (.A0(_1676_),
    .A1(\tms1x00.RAM[5][1] ),
    .S(_1718_),
    .X(_1720_));
 sky130_fd_sc_hd__clkbuf_1 _3678_ (.A(_1720_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _3679_ (.A0(_1678_),
    .A1(\tms1x00.RAM[5][2] ),
    .S(_1718_),
    .X(_1721_));
 sky130_fd_sc_hd__clkbuf_1 _3680_ (.A(_1721_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _3681_ (.A0(_1680_),
    .A1(\tms1x00.RAM[5][3] ),
    .S(_1718_),
    .X(_1722_));
 sky130_fd_sc_hd__clkbuf_1 _3682_ (.A(_1722_),
    .X(_0378_));
 sky130_fd_sc_hd__nor2_2 _3683_ (.A(_1233_),
    .B(_1263_),
    .Y(_1723_));
 sky130_fd_sc_hd__mux2_1 _3684_ (.A0(\tms1x00.RAM[67][0] ),
    .A1(_1629_),
    .S(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__clkbuf_1 _3685_ (.A(_1724_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _3686_ (.A0(\tms1x00.RAM[67][1] ),
    .A1(_1632_),
    .S(_1723_),
    .X(_1725_));
 sky130_fd_sc_hd__clkbuf_1 _3687_ (.A(_1725_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _3688_ (.A0(\tms1x00.RAM[67][2] ),
    .A1(_1634_),
    .S(_1723_),
    .X(_1726_));
 sky130_fd_sc_hd__clkbuf_1 _3689_ (.A(_1726_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _3690_ (.A0(\tms1x00.RAM[67][3] ),
    .A1(_1636_),
    .S(_1723_),
    .X(_1727_));
 sky130_fd_sc_hd__clkbuf_1 _3691_ (.A(_1727_),
    .X(_0382_));
 sky130_fd_sc_hd__or2_2 _3692_ (.A(_1263_),
    .B(_1271_),
    .X(_1728_));
 sky130_fd_sc_hd__mux2_1 _3693_ (.A0(_1673_),
    .A1(\tms1x00.RAM[66][0] ),
    .S(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__clkbuf_1 _3694_ (.A(_1729_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _3695_ (.A0(_1676_),
    .A1(\tms1x00.RAM[66][1] ),
    .S(_1728_),
    .X(_1730_));
 sky130_fd_sc_hd__clkbuf_1 _3696_ (.A(_1730_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _3697_ (.A0(_1678_),
    .A1(\tms1x00.RAM[66][2] ),
    .S(_1728_),
    .X(_1731_));
 sky130_fd_sc_hd__clkbuf_1 _3698_ (.A(_1731_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _3699_ (.A0(_1680_),
    .A1(\tms1x00.RAM[66][3] ),
    .S(_1728_),
    .X(_1732_));
 sky130_fd_sc_hd__clkbuf_1 _3700_ (.A(_1732_),
    .X(_0386_));
 sky130_fd_sc_hd__or4_4 _3701_ (.A(_0730_),
    .B(_0734_),
    .C(_0923_),
    .D(_1264_),
    .X(_1733_));
 sky130_fd_sc_hd__mux2_1 _3702_ (.A0(_1673_),
    .A1(\tms1x00.RAM[65][0] ),
    .S(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__clkbuf_1 _3703_ (.A(_1734_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _3704_ (.A0(_1676_),
    .A1(\tms1x00.RAM[65][1] ),
    .S(_1733_),
    .X(_1735_));
 sky130_fd_sc_hd__clkbuf_1 _3705_ (.A(_1735_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _3706_ (.A0(_1678_),
    .A1(\tms1x00.RAM[65][2] ),
    .S(_1733_),
    .X(_1736_));
 sky130_fd_sc_hd__clkbuf_1 _3707_ (.A(_1736_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _3708_ (.A0(_1680_),
    .A1(\tms1x00.RAM[65][3] ),
    .S(_1733_),
    .X(_1737_));
 sky130_fd_sc_hd__clkbuf_1 _3709_ (.A(_1737_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_2 _3710_ (.A(_1264_),
    .B(_1353_),
    .X(_1738_));
 sky130_fd_sc_hd__mux2_1 _3711_ (.A0(_1673_),
    .A1(\tms1x00.RAM[64][0] ),
    .S(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__clkbuf_1 _3712_ (.A(_1739_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _3713_ (.A0(_1676_),
    .A1(\tms1x00.RAM[64][1] ),
    .S(_1738_),
    .X(_1740_));
 sky130_fd_sc_hd__clkbuf_1 _3714_ (.A(_1740_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _3715_ (.A0(_1678_),
    .A1(\tms1x00.RAM[64][2] ),
    .S(_1738_),
    .X(_1741_));
 sky130_fd_sc_hd__clkbuf_1 _3716_ (.A(_1741_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _3717_ (.A0(_1680_),
    .A1(\tms1x00.RAM[64][3] ),
    .S(_1738_),
    .X(_1742_));
 sky130_fd_sc_hd__clkbuf_1 _3718_ (.A(_1742_),
    .X(_0394_));
 sky130_fd_sc_hd__or2_2 _3719_ (.A(_1284_),
    .B(_1403_),
    .X(_1743_));
 sky130_fd_sc_hd__mux2_1 _3720_ (.A0(_1673_),
    .A1(\tms1x00.RAM[63][0] ),
    .S(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__clkbuf_1 _3721_ (.A(_1744_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _3722_ (.A0(_1676_),
    .A1(\tms1x00.RAM[63][1] ),
    .S(_1743_),
    .X(_1745_));
 sky130_fd_sc_hd__clkbuf_1 _3723_ (.A(_1745_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _3724_ (.A0(_1678_),
    .A1(\tms1x00.RAM[63][2] ),
    .S(_1743_),
    .X(_1746_));
 sky130_fd_sc_hd__clkbuf_1 _3725_ (.A(_1746_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _3726_ (.A0(_1680_),
    .A1(\tms1x00.RAM[63][3] ),
    .S(_1743_),
    .X(_1747_));
 sky130_fd_sc_hd__clkbuf_1 _3727_ (.A(_1747_),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_4 _3728_ (.A(_0919_),
    .X(_1748_));
 sky130_fd_sc_hd__nor2_2 _3729_ (.A(_1264_),
    .B(_1316_),
    .Y(_1749_));
 sky130_fd_sc_hd__mux2_1 _3730_ (.A0(\tms1x00.RAM[71][0] ),
    .A1(_1748_),
    .S(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__clkbuf_1 _3731_ (.A(_1750_),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_4 _3732_ (.A(_1031_),
    .X(_1751_));
 sky130_fd_sc_hd__mux2_1 _3733_ (.A0(\tms1x00.RAM[71][1] ),
    .A1(_1751_),
    .S(_1749_),
    .X(_1752_));
 sky130_fd_sc_hd__clkbuf_1 _3734_ (.A(_1752_),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_4 _3735_ (.A(_1132_),
    .X(_1753_));
 sky130_fd_sc_hd__mux2_1 _3736_ (.A0(\tms1x00.RAM[71][2] ),
    .A1(_1753_),
    .S(_1749_),
    .X(_1754_));
 sky130_fd_sc_hd__clkbuf_1 _3737_ (.A(_1754_),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_4 _3738_ (.A(_1228_),
    .X(_1755_));
 sky130_fd_sc_hd__mux2_1 _3739_ (.A0(\tms1x00.RAM[71][3] ),
    .A1(_1755_),
    .S(_1749_),
    .X(_1756_));
 sky130_fd_sc_hd__clkbuf_1 _3740_ (.A(_1756_),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_4 _3741_ (.A(_0919_),
    .X(_1757_));
 sky130_fd_sc_hd__or2_2 _3742_ (.A(_1264_),
    .B(_1322_),
    .X(_1758_));
 sky130_fd_sc_hd__mux2_1 _3743_ (.A0(_1757_),
    .A1(\tms1x00.RAM[70][0] ),
    .S(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__clkbuf_1 _3744_ (.A(_1759_),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_4 _3745_ (.A(_1031_),
    .X(_1760_));
 sky130_fd_sc_hd__mux2_1 _3746_ (.A0(_1760_),
    .A1(\tms1x00.RAM[70][1] ),
    .S(_1758_),
    .X(_1761_));
 sky130_fd_sc_hd__clkbuf_1 _3747_ (.A(_1761_),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_4 _3748_ (.A(_1132_),
    .X(_1762_));
 sky130_fd_sc_hd__mux2_1 _3749_ (.A0(_1762_),
    .A1(\tms1x00.RAM[70][2] ),
    .S(_1758_),
    .X(_1763_));
 sky130_fd_sc_hd__clkbuf_1 _3750_ (.A(_1763_),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_4 _3751_ (.A(_1228_),
    .X(_1764_));
 sky130_fd_sc_hd__mux2_1 _3752_ (.A0(_1764_),
    .A1(\tms1x00.RAM[70][3] ),
    .S(_1758_),
    .X(_1765_));
 sky130_fd_sc_hd__clkbuf_1 _3753_ (.A(_1765_),
    .X(_0406_));
 sky130_fd_sc_hd__nor2_2 _3754_ (.A(_1322_),
    .B(_1473_),
    .Y(_1766_));
 sky130_fd_sc_hd__mux2_1 _3755_ (.A0(\tms1x00.RAM[6][0] ),
    .A1(_1748_),
    .S(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__clkbuf_1 _3756_ (.A(_1767_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _3757_ (.A0(\tms1x00.RAM[6][1] ),
    .A1(_1751_),
    .S(_1766_),
    .X(_1768_));
 sky130_fd_sc_hd__clkbuf_1 _3758_ (.A(_1768_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _3759_ (.A0(\tms1x00.RAM[6][2] ),
    .A1(_1753_),
    .S(_1766_),
    .X(_1769_));
 sky130_fd_sc_hd__clkbuf_1 _3760_ (.A(_1769_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _3761_ (.A0(\tms1x00.RAM[6][3] ),
    .A1(_1755_),
    .S(_1766_),
    .X(_1770_));
 sky130_fd_sc_hd__clkbuf_1 _3762_ (.A(_1770_),
    .X(_0410_));
 sky130_fd_sc_hd__or2_2 _3763_ (.A(_1264_),
    .B(_1337_),
    .X(_1771_));
 sky130_fd_sc_hd__mux2_1 _3764_ (.A0(_1757_),
    .A1(\tms1x00.RAM[68][0] ),
    .S(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__clkbuf_1 _3765_ (.A(_1772_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _3766_ (.A0(_1760_),
    .A1(\tms1x00.RAM[68][1] ),
    .S(_1771_),
    .X(_1773_));
 sky130_fd_sc_hd__clkbuf_1 _3767_ (.A(_1773_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _3768_ (.A0(_1762_),
    .A1(\tms1x00.RAM[68][2] ),
    .S(_1771_),
    .X(_1774_));
 sky130_fd_sc_hd__clkbuf_1 _3769_ (.A(_1774_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3770_ (.A0(_1764_),
    .A1(\tms1x00.RAM[68][3] ),
    .S(_1771_),
    .X(_1775_));
 sky130_fd_sc_hd__clkbuf_1 _3771_ (.A(_1775_),
    .X(_0414_));
 sky130_fd_sc_hd__or2_2 _3772_ (.A(_1263_),
    .B(_1422_),
    .X(_1776_));
 sky130_fd_sc_hd__mux2_1 _3773_ (.A0(_1757_),
    .A1(\tms1x00.RAM[76][0] ),
    .S(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__clkbuf_1 _3774_ (.A(_1777_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _3775_ (.A0(_1760_),
    .A1(\tms1x00.RAM[76][1] ),
    .S(_1776_),
    .X(_1778_));
 sky130_fd_sc_hd__clkbuf_1 _3776_ (.A(_1778_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _3777_ (.A0(_1762_),
    .A1(\tms1x00.RAM[76][2] ),
    .S(_1776_),
    .X(_1779_));
 sky130_fd_sc_hd__clkbuf_1 _3778_ (.A(_1779_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3779_ (.A0(_1764_),
    .A1(\tms1x00.RAM[76][3] ),
    .S(_1776_),
    .X(_1780_));
 sky130_fd_sc_hd__clkbuf_1 _3780_ (.A(_1780_),
    .X(_0418_));
 sky130_fd_sc_hd__nor2_2 _3781_ (.A(_1264_),
    .B(_1287_),
    .Y(_1781_));
 sky130_fd_sc_hd__mux2_1 _3782_ (.A0(\tms1x00.RAM[75][0] ),
    .A1(_1748_),
    .S(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__clkbuf_1 _3783_ (.A(_1782_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _3784_ (.A0(\tms1x00.RAM[75][1] ),
    .A1(_1751_),
    .S(_1781_),
    .X(_1783_));
 sky130_fd_sc_hd__clkbuf_1 _3785_ (.A(_1783_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _3786_ (.A0(\tms1x00.RAM[75][2] ),
    .A1(_1753_),
    .S(_1781_),
    .X(_1784_));
 sky130_fd_sc_hd__clkbuf_1 _3787_ (.A(_1784_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _3788_ (.A0(\tms1x00.RAM[75][3] ),
    .A1(_1755_),
    .S(_1781_),
    .X(_1785_));
 sky130_fd_sc_hd__clkbuf_1 _3789_ (.A(_1785_),
    .X(_0422_));
 sky130_fd_sc_hd__or2_2 _3790_ (.A(_1263_),
    .B(_1416_),
    .X(_1786_));
 sky130_fd_sc_hd__mux2_1 _3791_ (.A0(_1757_),
    .A1(\tms1x00.RAM[74][0] ),
    .S(_1786_),
    .X(_1787_));
 sky130_fd_sc_hd__clkbuf_1 _3792_ (.A(_1787_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _3793_ (.A0(_1760_),
    .A1(\tms1x00.RAM[74][1] ),
    .S(_1786_),
    .X(_1788_));
 sky130_fd_sc_hd__clkbuf_1 _3794_ (.A(_1788_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _3795_ (.A0(_1762_),
    .A1(\tms1x00.RAM[74][2] ),
    .S(_1786_),
    .X(_1789_));
 sky130_fd_sc_hd__clkbuf_1 _3796_ (.A(_1789_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _3797_ (.A0(_1764_),
    .A1(\tms1x00.RAM[74][3] ),
    .S(_1786_),
    .X(_1790_));
 sky130_fd_sc_hd__clkbuf_1 _3798_ (.A(_1790_),
    .X(_0426_));
 sky130_fd_sc_hd__or2_2 _3799_ (.A(_1255_),
    .B(_1263_),
    .X(_1791_));
 sky130_fd_sc_hd__mux2_1 _3800_ (.A0(_1757_),
    .A1(\tms1x00.RAM[73][0] ),
    .S(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__clkbuf_1 _3801_ (.A(_1792_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _3802_ (.A0(_1760_),
    .A1(\tms1x00.RAM[73][1] ),
    .S(_1791_),
    .X(_1793_));
 sky130_fd_sc_hd__clkbuf_1 _3803_ (.A(_1793_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _3804_ (.A0(_1762_),
    .A1(\tms1x00.RAM[73][2] ),
    .S(_1791_),
    .X(_1794_));
 sky130_fd_sc_hd__clkbuf_1 _3805_ (.A(_1794_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _3806_ (.A0(_1764_),
    .A1(\tms1x00.RAM[73][3] ),
    .S(_1791_),
    .X(_1795_));
 sky130_fd_sc_hd__clkbuf_1 _3807_ (.A(_1795_),
    .X(_0430_));
 sky130_fd_sc_hd__or2_2 _3808_ (.A(_1264_),
    .B(_1308_),
    .X(_1796_));
 sky130_fd_sc_hd__mux2_1 _3809_ (.A0(_1757_),
    .A1(\tms1x00.RAM[72][0] ),
    .S(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__clkbuf_1 _3810_ (.A(_1797_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _3811_ (.A0(_1760_),
    .A1(\tms1x00.RAM[72][1] ),
    .S(_1796_),
    .X(_1798_));
 sky130_fd_sc_hd__clkbuf_1 _3812_ (.A(_1798_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _3813_ (.A0(_1762_),
    .A1(\tms1x00.RAM[72][2] ),
    .S(_1796_),
    .X(_1799_));
 sky130_fd_sc_hd__clkbuf_1 _3814_ (.A(_1799_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _3815_ (.A0(_1764_),
    .A1(\tms1x00.RAM[72][3] ),
    .S(_1796_),
    .X(_1800_));
 sky130_fd_sc_hd__clkbuf_1 _3816_ (.A(_1800_),
    .X(_0434_));
 sky130_fd_sc_hd__nor2_2 _3817_ (.A(_1253_),
    .B(_1355_),
    .Y(_1801_));
 sky130_fd_sc_hd__mux2_1 _3818_ (.A0(\tms1x00.RAM[80][0] ),
    .A1(_1748_),
    .S(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__clkbuf_1 _3819_ (.A(_1802_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _3820_ (.A0(\tms1x00.RAM[80][1] ),
    .A1(_1751_),
    .S(_1801_),
    .X(_1803_));
 sky130_fd_sc_hd__clkbuf_1 _3821_ (.A(_1803_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _3822_ (.A0(\tms1x00.RAM[80][2] ),
    .A1(_1753_),
    .S(_1801_),
    .X(_1804_));
 sky130_fd_sc_hd__clkbuf_1 _3823_ (.A(_1804_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _3824_ (.A0(\tms1x00.RAM[80][3] ),
    .A1(_1755_),
    .S(_1801_),
    .X(_1805_));
 sky130_fd_sc_hd__clkbuf_1 _3825_ (.A(_1805_),
    .X(_0438_));
 sky130_fd_sc_hd__nor2_2 _3826_ (.A(_1316_),
    .B(_1473_),
    .Y(_1806_));
 sky130_fd_sc_hd__mux2_1 _3827_ (.A0(\tms1x00.RAM[7][0] ),
    .A1(_1748_),
    .S(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__clkbuf_1 _3828_ (.A(_1807_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _3829_ (.A0(\tms1x00.RAM[7][1] ),
    .A1(_1751_),
    .S(_1806_),
    .X(_1808_));
 sky130_fd_sc_hd__clkbuf_1 _3830_ (.A(_1808_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _3831_ (.A0(\tms1x00.RAM[7][2] ),
    .A1(_1753_),
    .S(_1806_),
    .X(_1809_));
 sky130_fd_sc_hd__clkbuf_1 _3832_ (.A(_1809_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _3833_ (.A0(\tms1x00.RAM[7][3] ),
    .A1(_1755_),
    .S(_1806_),
    .X(_1810_));
 sky130_fd_sc_hd__clkbuf_1 _3834_ (.A(_1810_),
    .X(_0442_));
 sky130_fd_sc_hd__or2_2 _3835_ (.A(_1263_),
    .B(_1410_),
    .X(_1811_));
 sky130_fd_sc_hd__mux2_1 _3836_ (.A0(_1757_),
    .A1(\tms1x00.RAM[78][0] ),
    .S(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__clkbuf_1 _3837_ (.A(_1812_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _3838_ (.A0(_1760_),
    .A1(\tms1x00.RAM[78][1] ),
    .S(_1811_),
    .X(_1813_));
 sky130_fd_sc_hd__clkbuf_1 _3839_ (.A(_1813_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _3840_ (.A0(_1762_),
    .A1(\tms1x00.RAM[78][2] ),
    .S(_1811_),
    .X(_1814_));
 sky130_fd_sc_hd__clkbuf_1 _3841_ (.A(_1814_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _3842_ (.A0(_1764_),
    .A1(\tms1x00.RAM[78][3] ),
    .S(_1811_),
    .X(_1815_));
 sky130_fd_sc_hd__clkbuf_1 _3843_ (.A(_1815_),
    .X(_0446_));
 sky130_fd_sc_hd__nor2_2 _3844_ (.A(_0928_),
    .B(_1263_),
    .Y(_1816_));
 sky130_fd_sc_hd__mux2_1 _3845_ (.A0(\tms1x00.RAM[77][0] ),
    .A1(_1748_),
    .S(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__clkbuf_1 _3846_ (.A(_1817_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _3847_ (.A0(\tms1x00.RAM[77][1] ),
    .A1(_1751_),
    .S(_1816_),
    .X(_1818_));
 sky130_fd_sc_hd__clkbuf_1 _3848_ (.A(_1818_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _3849_ (.A0(\tms1x00.RAM[77][2] ),
    .A1(_1753_),
    .S(_1816_),
    .X(_1819_));
 sky130_fd_sc_hd__clkbuf_1 _3850_ (.A(_1819_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _3851_ (.A0(\tms1x00.RAM[77][3] ),
    .A1(_1755_),
    .S(_1816_),
    .X(_1820_));
 sky130_fd_sc_hd__clkbuf_1 _3852_ (.A(_1820_),
    .X(_0450_));
 sky130_fd_sc_hd__or2_2 _3853_ (.A(_1253_),
    .B(_1278_),
    .X(_1821_));
 sky130_fd_sc_hd__mux2_1 _3854_ (.A0(_1757_),
    .A1(\tms1x00.RAM[85][0] ),
    .S(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__clkbuf_1 _3855_ (.A(_1822_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _3856_ (.A0(_1760_),
    .A1(\tms1x00.RAM[85][1] ),
    .S(_1821_),
    .X(_1823_));
 sky130_fd_sc_hd__clkbuf_1 _3857_ (.A(_1823_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _3858_ (.A0(_1762_),
    .A1(\tms1x00.RAM[85][2] ),
    .S(_1821_),
    .X(_1824_));
 sky130_fd_sc_hd__clkbuf_1 _3859_ (.A(_1824_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _3860_ (.A0(_1764_),
    .A1(\tms1x00.RAM[85][3] ),
    .S(_1821_),
    .X(_1825_));
 sky130_fd_sc_hd__clkbuf_1 _3861_ (.A(_1825_),
    .X(_0454_));
 sky130_fd_sc_hd__nor2_2 _3862_ (.A(_1253_),
    .B(_1339_),
    .Y(_1826_));
 sky130_fd_sc_hd__mux2_1 _3863_ (.A0(\tms1x00.RAM[84][0] ),
    .A1(_1748_),
    .S(_1826_),
    .X(_1827_));
 sky130_fd_sc_hd__clkbuf_1 _3864_ (.A(_1827_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _3865_ (.A0(\tms1x00.RAM[84][1] ),
    .A1(_1751_),
    .S(_1826_),
    .X(_1828_));
 sky130_fd_sc_hd__clkbuf_1 _3866_ (.A(_1828_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _3867_ (.A0(\tms1x00.RAM[84][2] ),
    .A1(_1753_),
    .S(_1826_),
    .X(_1829_));
 sky130_fd_sc_hd__clkbuf_1 _3868_ (.A(_1829_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _3869_ (.A0(\tms1x00.RAM[84][3] ),
    .A1(_1755_),
    .S(_1826_),
    .X(_1830_));
 sky130_fd_sc_hd__clkbuf_1 _3870_ (.A(_1830_),
    .X(_0458_));
 sky130_fd_sc_hd__nor2_2 _3871_ (.A(_1233_),
    .B(_1253_),
    .Y(_1831_));
 sky130_fd_sc_hd__mux2_1 _3872_ (.A0(\tms1x00.RAM[83][0] ),
    .A1(_1748_),
    .S(_1831_),
    .X(_1832_));
 sky130_fd_sc_hd__clkbuf_1 _3873_ (.A(_1832_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _3874_ (.A0(\tms1x00.RAM[83][1] ),
    .A1(_1751_),
    .S(_1831_),
    .X(_1833_));
 sky130_fd_sc_hd__clkbuf_1 _3875_ (.A(_1833_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _3876_ (.A0(\tms1x00.RAM[83][2] ),
    .A1(_1753_),
    .S(_1831_),
    .X(_1834_));
 sky130_fd_sc_hd__clkbuf_1 _3877_ (.A(_1834_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _3878_ (.A0(\tms1x00.RAM[83][3] ),
    .A1(_1755_),
    .S(_1831_),
    .X(_1835_));
 sky130_fd_sc_hd__clkbuf_1 _3879_ (.A(_1835_),
    .X(_0462_));
 sky130_fd_sc_hd__or2_2 _3880_ (.A(_1253_),
    .B(_1271_),
    .X(_1836_));
 sky130_fd_sc_hd__mux2_1 _3881_ (.A0(_1757_),
    .A1(\tms1x00.RAM[82][0] ),
    .S(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__clkbuf_1 _3882_ (.A(_1837_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _3883_ (.A0(_1760_),
    .A1(\tms1x00.RAM[82][1] ),
    .S(_1836_),
    .X(_1838_));
 sky130_fd_sc_hd__clkbuf_1 _3884_ (.A(_1838_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _3885_ (.A0(_1762_),
    .A1(\tms1x00.RAM[82][2] ),
    .S(_1836_),
    .X(_1839_));
 sky130_fd_sc_hd__clkbuf_1 _3886_ (.A(_1839_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _3887_ (.A0(_1764_),
    .A1(\tms1x00.RAM[82][3] ),
    .S(_1836_),
    .X(_1840_));
 sky130_fd_sc_hd__clkbuf_1 _3888_ (.A(_1840_),
    .X(_0466_));
 sky130_fd_sc_hd__or2_2 _3889_ (.A(_1286_),
    .B(_1252_),
    .X(_1841_));
 sky130_fd_sc_hd__nor4_4 _3890_ (.A(_0730_),
    .B(_0734_),
    .C(_0923_),
    .D(_1841_),
    .Y(_1842_));
 sky130_fd_sc_hd__mux2_1 _3891_ (.A0(\tms1x00.RAM[81][0] ),
    .A1(_1748_),
    .S(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__clkbuf_1 _3892_ (.A(_1843_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _3893_ (.A0(\tms1x00.RAM[81][1] ),
    .A1(_1751_),
    .S(_1842_),
    .X(_1844_));
 sky130_fd_sc_hd__clkbuf_1 _3894_ (.A(_1844_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _3895_ (.A0(\tms1x00.RAM[81][2] ),
    .A1(_1753_),
    .S(_1842_),
    .X(_1845_));
 sky130_fd_sc_hd__clkbuf_1 _3896_ (.A(_1845_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _3897_ (.A0(\tms1x00.RAM[81][3] ),
    .A1(_1755_),
    .S(_1842_),
    .X(_1846_));
 sky130_fd_sc_hd__clkbuf_1 _3898_ (.A(_1846_),
    .X(_0470_));
 sky130_fd_sc_hd__nor2_2 _3899_ (.A(_1253_),
    .B(_1324_),
    .Y(_1847_));
 sky130_fd_sc_hd__mux2_1 _3900_ (.A0(\tms1x00.RAM[86][0] ),
    .A1(_1748_),
    .S(_1847_),
    .X(_1848_));
 sky130_fd_sc_hd__clkbuf_1 _3901_ (.A(_1848_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _3902_ (.A0(\tms1x00.RAM[86][1] ),
    .A1(_1751_),
    .S(_1847_),
    .X(_1849_));
 sky130_fd_sc_hd__clkbuf_1 _3903_ (.A(_1849_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _3904_ (.A0(\tms1x00.RAM[86][2] ),
    .A1(_1753_),
    .S(_1847_),
    .X(_1850_));
 sky130_fd_sc_hd__clkbuf_1 _3905_ (.A(_1850_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _3906_ (.A0(\tms1x00.RAM[86][3] ),
    .A1(_1755_),
    .S(_1847_),
    .X(_1851_));
 sky130_fd_sc_hd__clkbuf_1 _3907_ (.A(_1851_),
    .X(_0474_));
 sky130_fd_sc_hd__nor2_2 _3908_ (.A(_1308_),
    .B(_1473_),
    .Y(_1852_));
 sky130_fd_sc_hd__mux2_1 _3909_ (.A0(\tms1x00.RAM[8][0] ),
    .A1(_1335_),
    .S(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__clkbuf_1 _3910_ (.A(_1853_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _3911_ (.A0(\tms1x00.RAM[8][1] ),
    .A1(_1342_),
    .S(_1852_),
    .X(_1854_));
 sky130_fd_sc_hd__clkbuf_1 _3912_ (.A(_1854_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _3913_ (.A0(\tms1x00.RAM[8][2] ),
    .A1(_1345_),
    .S(_1852_),
    .X(_1855_));
 sky130_fd_sc_hd__clkbuf_1 _3914_ (.A(_1855_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _3915_ (.A0(\tms1x00.RAM[8][3] ),
    .A1(_1348_),
    .S(_1852_),
    .X(_1856_));
 sky130_fd_sc_hd__clkbuf_1 _3916_ (.A(_1856_),
    .X(_0478_));
 sky130_fd_sc_hd__or2_2 _3917_ (.A(_1253_),
    .B(_1309_),
    .X(_1857_));
 sky130_fd_sc_hd__mux2_1 _3918_ (.A0(_1757_),
    .A1(\tms1x00.RAM[88][0] ),
    .S(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__clkbuf_1 _3919_ (.A(_1858_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _3920_ (.A0(_1760_),
    .A1(\tms1x00.RAM[88][1] ),
    .S(_1857_),
    .X(_1859_));
 sky130_fd_sc_hd__clkbuf_1 _3921_ (.A(_1859_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _3922_ (.A0(_1762_),
    .A1(\tms1x00.RAM[88][2] ),
    .S(_1857_),
    .X(_1860_));
 sky130_fd_sc_hd__clkbuf_1 _3923_ (.A(_1860_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _3924_ (.A0(_1764_),
    .A1(\tms1x00.RAM[88][3] ),
    .S(_1857_),
    .X(_1861_));
 sky130_fd_sc_hd__clkbuf_1 _3925_ (.A(_1861_),
    .X(_0482_));
 sky130_fd_sc_hd__nor2_2 _3926_ (.A(_1316_),
    .B(_1841_),
    .Y(_1862_));
 sky130_fd_sc_hd__mux2_1 _3927_ (.A0(\tms1x00.RAM[87][0] ),
    .A1(_1335_),
    .S(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__clkbuf_1 _3928_ (.A(_1863_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _3929_ (.A0(\tms1x00.RAM[87][1] ),
    .A1(_1342_),
    .S(_1862_),
    .X(_1864_));
 sky130_fd_sc_hd__clkbuf_1 _3930_ (.A(_1864_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _3931_ (.A0(\tms1x00.RAM[87][2] ),
    .A1(_1345_),
    .S(_1862_),
    .X(_1865_));
 sky130_fd_sc_hd__clkbuf_1 _3932_ (.A(_1865_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _3933_ (.A0(\tms1x00.RAM[87][3] ),
    .A1(_1348_),
    .S(_1862_),
    .X(_1866_));
 sky130_fd_sc_hd__clkbuf_1 _3934_ (.A(_1866_),
    .X(_0486_));
 sky130_fd_sc_hd__buf_2 _3935_ (.A(_0919_),
    .X(_1867_));
 sky130_fd_sc_hd__or2_2 _3936_ (.A(_1252_),
    .B(_1410_),
    .X(_1868_));
 sky130_fd_sc_hd__mux2_1 _3937_ (.A0(_1867_),
    .A1(\tms1x00.RAM[94][0] ),
    .S(_1868_),
    .X(_1869_));
 sky130_fd_sc_hd__clkbuf_1 _3938_ (.A(_1869_),
    .X(_0487_));
 sky130_fd_sc_hd__buf_2 _3939_ (.A(_1031_),
    .X(_1870_));
 sky130_fd_sc_hd__mux2_1 _3940_ (.A0(_1870_),
    .A1(\tms1x00.RAM[94][1] ),
    .S(_1868_),
    .X(_1871_));
 sky130_fd_sc_hd__clkbuf_1 _3941_ (.A(_1871_),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_4 _3942_ (.A(_1132_),
    .X(_1872_));
 sky130_fd_sc_hd__mux2_1 _3943_ (.A0(_1872_),
    .A1(\tms1x00.RAM[94][2] ),
    .S(_1868_),
    .X(_1873_));
 sky130_fd_sc_hd__clkbuf_1 _3944_ (.A(_1873_),
    .X(_0489_));
 sky130_fd_sc_hd__clkbuf_4 _3945_ (.A(_1228_),
    .X(_1874_));
 sky130_fd_sc_hd__mux2_1 _3946_ (.A0(_1874_),
    .A1(\tms1x00.RAM[94][3] ),
    .S(_1868_),
    .X(_1875_));
 sky130_fd_sc_hd__clkbuf_1 _3947_ (.A(_1875_),
    .X(_0490_));
 sky130_fd_sc_hd__nor2_2 _3948_ (.A(_0928_),
    .B(_1253_),
    .Y(_1876_));
 sky130_fd_sc_hd__mux2_1 _3949_ (.A0(\tms1x00.RAM[93][0] ),
    .A1(_1335_),
    .S(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__clkbuf_1 _3950_ (.A(_1877_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _3951_ (.A0(\tms1x00.RAM[93][1] ),
    .A1(_1342_),
    .S(_1876_),
    .X(_1878_));
 sky130_fd_sc_hd__clkbuf_1 _3952_ (.A(_1878_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _3953_ (.A0(\tms1x00.RAM[93][2] ),
    .A1(_1345_),
    .S(_1876_),
    .X(_1879_));
 sky130_fd_sc_hd__clkbuf_1 _3954_ (.A(_1879_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _3955_ (.A0(\tms1x00.RAM[93][3] ),
    .A1(_1348_),
    .S(_1876_),
    .X(_1880_));
 sky130_fd_sc_hd__clkbuf_1 _3956_ (.A(_1880_),
    .X(_0494_));
 sky130_fd_sc_hd__or2_2 _3957_ (.A(_1252_),
    .B(_1422_),
    .X(_1881_));
 sky130_fd_sc_hd__mux2_1 _3958_ (.A0(_1867_),
    .A1(\tms1x00.RAM[92][0] ),
    .S(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__clkbuf_1 _3959_ (.A(_1882_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _3960_ (.A0(_1870_),
    .A1(\tms1x00.RAM[92][1] ),
    .S(_1881_),
    .X(_1883_));
 sky130_fd_sc_hd__clkbuf_1 _3961_ (.A(_1883_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _3962_ (.A0(_1872_),
    .A1(\tms1x00.RAM[92][2] ),
    .S(_1881_),
    .X(_1884_));
 sky130_fd_sc_hd__clkbuf_1 _3963_ (.A(_1884_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _3964_ (.A0(_1874_),
    .A1(\tms1x00.RAM[92][3] ),
    .S(_1881_),
    .X(_1885_));
 sky130_fd_sc_hd__clkbuf_1 _3965_ (.A(_1885_),
    .X(_0498_));
 sky130_fd_sc_hd__or2_2 _3966_ (.A(_1252_),
    .B(_1288_),
    .X(_1886_));
 sky130_fd_sc_hd__mux2_1 _3967_ (.A0(_1867_),
    .A1(\tms1x00.RAM[91][0] ),
    .S(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__clkbuf_1 _3968_ (.A(_1887_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _3969_ (.A0(_1870_),
    .A1(\tms1x00.RAM[91][1] ),
    .S(_1886_),
    .X(_1888_));
 sky130_fd_sc_hd__clkbuf_1 _3970_ (.A(_1888_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _3971_ (.A0(_1872_),
    .A1(\tms1x00.RAM[91][2] ),
    .S(_1886_),
    .X(_1889_));
 sky130_fd_sc_hd__clkbuf_1 _3972_ (.A(_1889_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _3973_ (.A0(_1874_),
    .A1(\tms1x00.RAM[91][3] ),
    .S(_1886_),
    .X(_1890_));
 sky130_fd_sc_hd__clkbuf_1 _3974_ (.A(_1890_),
    .X(_0502_));
 sky130_fd_sc_hd__or2_2 _3975_ (.A(_1252_),
    .B(_1416_),
    .X(_1891_));
 sky130_fd_sc_hd__mux2_1 _3976_ (.A0(_1867_),
    .A1(\tms1x00.RAM[90][0] ),
    .S(_1891_),
    .X(_1892_));
 sky130_fd_sc_hd__clkbuf_1 _3977_ (.A(_1892_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _3978_ (.A0(_1870_),
    .A1(\tms1x00.RAM[90][1] ),
    .S(_1891_),
    .X(_1893_));
 sky130_fd_sc_hd__clkbuf_1 _3979_ (.A(_1893_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _3980_ (.A0(_1872_),
    .A1(\tms1x00.RAM[90][2] ),
    .S(_1891_),
    .X(_1894_));
 sky130_fd_sc_hd__clkbuf_1 _3981_ (.A(_1894_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _3982_ (.A0(_1874_),
    .A1(\tms1x00.RAM[90][3] ),
    .S(_1891_),
    .X(_1895_));
 sky130_fd_sc_hd__clkbuf_1 _3983_ (.A(_1895_),
    .X(_0506_));
 sky130_fd_sc_hd__or3_4 _3984_ (.A(_1286_),
    .B(_1240_),
    .C(_1316_),
    .X(_1896_));
 sky130_fd_sc_hd__mux2_1 _3985_ (.A0(_1867_),
    .A1(\tms1x00.RAM[23][0] ),
    .S(_1896_),
    .X(_1897_));
 sky130_fd_sc_hd__clkbuf_1 _3986_ (.A(_1897_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _3987_ (.A0(_1870_),
    .A1(\tms1x00.RAM[23][1] ),
    .S(_1896_),
    .X(_1898_));
 sky130_fd_sc_hd__clkbuf_1 _3988_ (.A(_1898_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _3989_ (.A0(_1872_),
    .A1(\tms1x00.RAM[23][2] ),
    .S(_1896_),
    .X(_1899_));
 sky130_fd_sc_hd__clkbuf_1 _3990_ (.A(_1899_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _3991_ (.A0(_1874_),
    .A1(\tms1x00.RAM[23][3] ),
    .S(_1896_),
    .X(_1900_));
 sky130_fd_sc_hd__clkbuf_1 _3992_ (.A(_1900_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _3993_ (.A0(\tms1x00.Y[0] ),
    .A1(_0720_),
    .S(_0725_),
    .X(_1901_));
 sky130_fd_sc_hd__clkbuf_1 _3994_ (.A(_1901_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _3995_ (.A0(\tms1x00.Y[1] ),
    .A1(_0727_),
    .S(_0725_),
    .X(_1902_));
 sky130_fd_sc_hd__clkbuf_1 _3996_ (.A(_1902_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _3997_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0725_),
    .X(_1903_));
 sky130_fd_sc_hd__clkbuf_1 _3998_ (.A(_1903_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _3999_ (.A0(_0733_),
    .A1(_0734_),
    .S(_0724_),
    .X(_1904_));
 sky130_fd_sc_hd__clkbuf_1 _4000_ (.A(_1904_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _4001_ (.A0(\tms1x00.X[2] ),
    .A1(\tms1x00.ram_addr_buff[4] ),
    .S(_0724_),
    .X(_1905_));
 sky130_fd_sc_hd__clkbuf_1 _4002_ (.A(_1905_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _4003_ (.A0(\tms1x00.X[0] ),
    .A1(\tms1x00.ram_addr_buff[5] ),
    .S(_0724_),
    .X(_1906_));
 sky130_fd_sc_hd__clkbuf_1 _4004_ (.A(_1906_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _4005_ (.A0(\tms1x00.X[1] ),
    .A1(\tms1x00.ram_addr_buff[6] ),
    .S(_0724_),
    .X(_1907_));
 sky130_fd_sc_hd__clkbuf_1 _4006_ (.A(_1907_),
    .X(_0517_));
 sky130_fd_sc_hd__and2_1 _4007_ (.A(\tms1x00.wb_step ),
    .B(_0762_),
    .X(_1908_));
 sky130_fd_sc_hd__clkbuf_1 _4008_ (.A(_1908_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _4009_ (.A0(net1),
    .A1(chip_sel_override),
    .S(net152),
    .X(_1909_));
 sky130_fd_sc_hd__buf_2 _4010_ (.A(_0719_),
    .X(_1910_));
 sky130_fd_sc_hd__mux2_1 _4011_ (.A0(net96),
    .A1(_1909_),
    .S(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__clkbuf_1 _4012_ (.A(_1911_),
    .X(_0519_));
 sky130_fd_sc_hd__mux4_1 _4013_ (.A0(net6),
    .A1(net8),
    .A2(net9),
    .A3(net10),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_1912_));
 sky130_fd_sc_hd__nor2_4 _4014_ (.A(_0721_),
    .B(_0745_),
    .Y(_1913_));
 sky130_fd_sc_hd__mux2_1 _4015_ (.A0(\tms1x00.ins_in[0] ),
    .A1(_1912_),
    .S(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__or2_1 _4016_ (.A(net106),
    .B(_1914_),
    .X(_1915_));
 sky130_fd_sc_hd__clkbuf_1 _4017_ (.A(_1915_),
    .X(_0520_));
 sky130_fd_sc_hd__mux4_1 _4018_ (.A0(net8),
    .A1(net9),
    .A2(net10),
    .A3(net11),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_1916_));
 sky130_fd_sc_hd__mux2_1 _4019_ (.A0(\tms1x00.ins_in[1] ),
    .A1(_1916_),
    .S(_1913_),
    .X(_1917_));
 sky130_fd_sc_hd__or2_1 _4020_ (.A(net106),
    .B(_1917_),
    .X(_1918_));
 sky130_fd_sc_hd__clkbuf_1 _4021_ (.A(_1918_),
    .X(_0521_));
 sky130_fd_sc_hd__or2_1 _4022_ (.A(_0721_),
    .B(_0745_),
    .X(_1919_));
 sky130_fd_sc_hd__mux4_1 _4023_ (.A0(net9),
    .A1(net10),
    .A2(net11),
    .A3(net12),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_1920_));
 sky130_fd_sc_hd__or2_1 _4024_ (.A(_1919_),
    .B(_1920_),
    .X(_1921_));
 sky130_fd_sc_hd__buf_2 _4025_ (.A(_0718_),
    .X(_1922_));
 sky130_fd_sc_hd__clkbuf_4 _4026_ (.A(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__o211a_1 _4027_ (.A1(\tms1x00.ins_in[2] ),
    .A2(_1913_),
    .B1(_1921_),
    .C1(_1923_),
    .X(_0522_));
 sky130_fd_sc_hd__mux4_1 _4028_ (.A0(net10),
    .A1(net11),
    .A2(net12),
    .A3(net13),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_1924_));
 sky130_fd_sc_hd__or2_1 _4029_ (.A(_1919_),
    .B(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__o211a_1 _4030_ (.A1(\tms1x00.ins_in[3] ),
    .A2(_1913_),
    .B1(_1925_),
    .C1(_1923_),
    .X(_0523_));
 sky130_fd_sc_hd__mux4_1 _4031_ (.A0(net11),
    .A1(net12),
    .A2(net13),
    .A3(net14),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_1926_));
 sky130_fd_sc_hd__or2_1 _4032_ (.A(_1919_),
    .B(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__o211a_1 _4033_ (.A1(_0743_),
    .A2(_1913_),
    .B1(_1927_),
    .C1(_1923_),
    .X(_0524_));
 sky130_fd_sc_hd__buf_2 _4034_ (.A(\tms1x00.ins_in[5] ),
    .X(_1928_));
 sky130_fd_sc_hd__mux4_1 _4035_ (.A0(net12),
    .A1(net13),
    .A2(net14),
    .A3(net15),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_1929_));
 sky130_fd_sc_hd__mux2_1 _4036_ (.A0(_1928_),
    .A1(_1929_),
    .S(_1913_),
    .X(_1930_));
 sky130_fd_sc_hd__or2_1 _4037_ (.A(net106),
    .B(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_1 _4038_ (.A(_1931_),
    .X(_0525_));
 sky130_fd_sc_hd__mux4_1 _4039_ (.A0(net13),
    .A1(net14),
    .A2(net15),
    .A3(net16),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_1932_));
 sky130_fd_sc_hd__or2_1 _4040_ (.A(_1919_),
    .B(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__o211a_1 _4041_ (.A1(\tms1x00.ins_in[6] ),
    .A2(_1913_),
    .B1(_1933_),
    .C1(_1923_),
    .X(_0526_));
 sky130_fd_sc_hd__mux4_1 _4042_ (.A0(net14),
    .A1(net15),
    .A2(net16),
    .A3(net7),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_1934_));
 sky130_fd_sc_hd__or2_1 _4043_ (.A(_1919_),
    .B(_1934_),
    .X(_1935_));
 sky130_fd_sc_hd__o211a_1 _4044_ (.A1(_0742_),
    .A2(_1913_),
    .B1(_1935_),
    .C1(_1923_),
    .X(_0527_));
 sky130_fd_sc_hd__nand2_2 _4045_ (.A(net152),
    .B(_0722_),
    .Y(_1936_));
 sky130_fd_sc_hd__nand2_1 _4046_ (.A(net151),
    .B(_1936_),
    .Y(_1937_));
 sky130_fd_sc_hd__or2_1 _4047_ (.A(net151),
    .B(_1936_),
    .X(_1938_));
 sky130_fd_sc_hd__and3_1 _4048_ (.A(_0762_),
    .B(_1937_),
    .C(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__clkbuf_1 _4049_ (.A(_1939_),
    .X(_0528_));
 sky130_fd_sc_hd__nor2_1 _4050_ (.A(net79),
    .B(net78),
    .Y(_1940_));
 sky130_fd_sc_hd__a21o_1 _4051_ (.A1(net151),
    .A2(_1936_),
    .B1(net78),
    .X(_1941_));
 sky130_fd_sc_hd__o211a_1 _4052_ (.A1(_1937_),
    .A2(_1940_),
    .B1(_1941_),
    .C1(_1923_),
    .X(_0529_));
 sky130_fd_sc_hd__a21oi_1 _4053_ (.A1(net79),
    .A2(_1937_),
    .B1(_0757_),
    .Y(_1942_));
 sky130_fd_sc_hd__nor2_1 _4054_ (.A(net106),
    .B(_1942_),
    .Y(_0530_));
 sky130_fd_sc_hd__and2b_1 _4055_ (.A_N(\tms1x00.Y[1] ),
    .B(\tms1x00.Y[0] ),
    .X(_1943_));
 sky130_fd_sc_hd__a41o_1 _4056_ (.A1(_0753_),
    .A2(_0739_),
    .A3(_0759_),
    .A4(_1943_),
    .B1(net81),
    .X(_1944_));
 sky130_fd_sc_hd__or4b_1 _4057_ (.A(_0732_),
    .B(_0729_),
    .C(_0750_),
    .D_N(_1943_),
    .X(_1945_));
 sky130_fd_sc_hd__and3_1 _4058_ (.A(_1922_),
    .B(_1944_),
    .C(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__clkbuf_1 _4059_ (.A(_1946_),
    .X(_0531_));
 sky130_fd_sc_hd__and2b_1 _4060_ (.A_N(\tms1x00.Y[0] ),
    .B(\tms1x00.Y[1] ),
    .X(_1947_));
 sky130_fd_sc_hd__a41o_1 _4061_ (.A1(_0752_),
    .A2(_0739_),
    .A3(_0759_),
    .A4(_1947_),
    .B1(net82),
    .X(_1948_));
 sky130_fd_sc_hd__or4b_1 _4062_ (.A(\tms1x00.Y[3] ),
    .B(_0729_),
    .C(_0750_),
    .D_N(_1947_),
    .X(_1949_));
 sky130_fd_sc_hd__and3_1 _4063_ (.A(_1922_),
    .B(_1948_),
    .C(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__clkbuf_1 _4064_ (.A(_1950_),
    .X(_0532_));
 sky130_fd_sc_hd__nand2_1 _4065_ (.A(\tms1x00.Y[1] ),
    .B(\tms1x00.Y[0] ),
    .Y(_1951_));
 sky130_fd_sc_hd__nor2_1 _4066_ (.A(\tms1x00.Y[2] ),
    .B(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__and2_1 _4067_ (.A(_0752_),
    .B(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__a21o_1 _4068_ (.A1(_0760_),
    .A2(_1953_),
    .B1(net83),
    .X(_1954_));
 sky130_fd_sc_hd__or2b_1 _4069_ (.A(_0751_),
    .B_N(_1953_),
    .X(_1955_));
 sky130_fd_sc_hd__and3_1 _4070_ (.A(_1922_),
    .B(_1954_),
    .C(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__clkbuf_1 _4071_ (.A(_1956_),
    .X(_0533_));
 sky130_fd_sc_hd__or3b_1 _4072_ (.A(_0732_),
    .B(_0739_),
    .C_N(_0740_),
    .X(_1957_));
 sky130_fd_sc_hd__a41o_1 _4073_ (.A1(_0753_),
    .A2(_0729_),
    .A3(_0740_),
    .A4(_0760_),
    .B1(net84),
    .X(_1958_));
 sky130_fd_sc_hd__o211a_1 _4074_ (.A1(_0751_),
    .A2(_1957_),
    .B1(_1958_),
    .C1(_1923_),
    .X(_0534_));
 sky130_fd_sc_hd__nand2_1 _4075_ (.A(\tms1x00.Y[2] ),
    .B(_1943_),
    .Y(_1959_));
 sky130_fd_sc_hd__inv_2 _4076_ (.A(_1959_),
    .Y(_1960_));
 sky130_fd_sc_hd__and3_1 _4077_ (.A(_0753_),
    .B(_0759_),
    .C(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__o21a_1 _4078_ (.A1(net85),
    .A2(_1961_),
    .B1(_0762_),
    .X(_1962_));
 sky130_fd_sc_hd__o31a_1 _4079_ (.A1(_0733_),
    .A2(_0751_),
    .A3(_1959_),
    .B1(_1962_),
    .X(_0535_));
 sky130_fd_sc_hd__nand2_1 _4080_ (.A(\tms1x00.Y[2] ),
    .B(_1947_),
    .Y(_1963_));
 sky130_fd_sc_hd__inv_2 _4081_ (.A(_1963_),
    .Y(_1964_));
 sky130_fd_sc_hd__and3_1 _4082_ (.A(_0753_),
    .B(_0759_),
    .C(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__o21a_1 _4083_ (.A1(net86),
    .A2(_1965_),
    .B1(_0762_),
    .X(_1966_));
 sky130_fd_sc_hd__o31a_1 _4084_ (.A1(_0733_),
    .A2(_0751_),
    .A3(_1963_),
    .B1(_1966_),
    .X(_0536_));
 sky130_fd_sc_hd__nor2_1 _4085_ (.A(_0739_),
    .B(_1951_),
    .Y(_1967_));
 sky130_fd_sc_hd__a31o_1 _4086_ (.A1(_0753_),
    .A2(_0760_),
    .A3(_1967_),
    .B1(net87),
    .X(_1968_));
 sky130_fd_sc_hd__or3b_1 _4087_ (.A(_0732_),
    .B(_0750_),
    .C_N(_1967_),
    .X(_1969_));
 sky130_fd_sc_hd__and3_1 _4088_ (.A(_1922_),
    .B(_1968_),
    .C(_1969_),
    .X(_1970_));
 sky130_fd_sc_hd__clkbuf_1 _4089_ (.A(_1970_),
    .X(_0537_));
 sky130_fd_sc_hd__a31o_1 _4090_ (.A1(_0733_),
    .A2(_0754_),
    .A3(_0760_),
    .B1(net88),
    .X(_1971_));
 sky130_fd_sc_hd__o311a_1 _4091_ (.A1(_0753_),
    .A2(_0741_),
    .A3(_0751_),
    .B1(_1971_),
    .C1(_0762_),
    .X(_0538_));
 sky130_fd_sc_hd__or3b_1 _4092_ (.A(_0753_),
    .B(_0729_),
    .C_N(_1943_),
    .X(_1972_));
 sky130_fd_sc_hd__a41o_1 _4093_ (.A1(_0733_),
    .A2(_0739_),
    .A3(_0760_),
    .A4(_1943_),
    .B1(net89),
    .X(_1973_));
 sky130_fd_sc_hd__o211a_1 _4094_ (.A1(_0751_),
    .A2(_1972_),
    .B1(_1973_),
    .C1(_1923_),
    .X(_0539_));
 sky130_fd_sc_hd__or3b_1 _4095_ (.A(_0753_),
    .B(_0729_),
    .C_N(_1947_),
    .X(_1974_));
 sky130_fd_sc_hd__a41o_1 _4096_ (.A1(_0732_),
    .A2(_0739_),
    .A3(_0760_),
    .A4(_1947_),
    .B1(net90),
    .X(_1975_));
 sky130_fd_sc_hd__o211a_1 _4097_ (.A1(_0751_),
    .A2(_1974_),
    .B1(_1975_),
    .C1(_1923_),
    .X(_0540_));
 sky130_fd_sc_hd__a31o_1 _4098_ (.A1(_0732_),
    .A2(_0760_),
    .A3(_1952_),
    .B1(net91),
    .X(_1976_));
 sky130_fd_sc_hd__or3b_1 _4099_ (.A(_0752_),
    .B(_0750_),
    .C_N(_1952_),
    .X(_1977_));
 sky130_fd_sc_hd__and3_1 _4100_ (.A(_1922_),
    .B(_1976_),
    .C(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__clkbuf_1 _4101_ (.A(_1978_),
    .X(_0541_));
 sky130_fd_sc_hd__or3b_1 _4102_ (.A(_0753_),
    .B(_0739_),
    .C_N(_0740_),
    .X(_1979_));
 sky130_fd_sc_hd__a41o_1 _4103_ (.A1(_0732_),
    .A2(_0729_),
    .A3(_0740_),
    .A4(_0760_),
    .B1(net92),
    .X(_1980_));
 sky130_fd_sc_hd__o211a_1 _4104_ (.A1(_0751_),
    .A2(_1979_),
    .B1(_1980_),
    .C1(_1923_),
    .X(_0542_));
 sky130_fd_sc_hd__a31o_1 _4105_ (.A1(_0732_),
    .A2(_0759_),
    .A3(_1960_),
    .B1(net93),
    .X(_1981_));
 sky130_fd_sc_hd__or3_1 _4106_ (.A(_0752_),
    .B(_0750_),
    .C(_1959_),
    .X(_1982_));
 sky130_fd_sc_hd__and3_1 _4107_ (.A(_1922_),
    .B(_1981_),
    .C(_1982_),
    .X(_1983_));
 sky130_fd_sc_hd__clkbuf_1 _4108_ (.A(_1983_),
    .X(_0543_));
 sky130_fd_sc_hd__a31o_1 _4109_ (.A1(_0732_),
    .A2(_0759_),
    .A3(_1964_),
    .B1(net94),
    .X(_1984_));
 sky130_fd_sc_hd__or3_1 _4110_ (.A(_0752_),
    .B(_0750_),
    .C(_1963_),
    .X(_1985_));
 sky130_fd_sc_hd__and3_1 _4111_ (.A(_1922_),
    .B(_1984_),
    .C(_1985_),
    .X(_1986_));
 sky130_fd_sc_hd__clkbuf_1 _4112_ (.A(_1986_),
    .X(_0544_));
 sky130_fd_sc_hd__nand2_1 _4113_ (.A(_0733_),
    .B(_1967_),
    .Y(_1987_));
 sky130_fd_sc_hd__a31o_1 _4114_ (.A1(_0733_),
    .A2(_0760_),
    .A3(_1967_),
    .B1(net95),
    .X(_1988_));
 sky130_fd_sc_hd__clkbuf_4 _4115_ (.A(_1922_),
    .X(_1989_));
 sky130_fd_sc_hd__o211a_1 _4116_ (.A1(_0751_),
    .A2(_1987_),
    .B1(_1988_),
    .C1(_1989_),
    .X(_0545_));
 sky130_fd_sc_hd__and2b_1 _4117_ (.A_N(_1928_),
    .B(_0743_),
    .X(_1990_));
 sky130_fd_sc_hd__nor3b_2 _4118_ (.A(_0763_),
    .B(_0749_),
    .C_N(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__or3b_2 _4119_ (.A(_0763_),
    .B(_0749_),
    .C_N(_1990_),
    .X(_1992_));
 sky130_fd_sc_hd__a21o_1 _4120_ (.A1(_0755_),
    .A2(\tms1x00.A[0] ),
    .B1(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__o211a_1 _4121_ (.A1(net72),
    .A2(_1991_),
    .B1(_1993_),
    .C1(_1989_),
    .X(_0546_));
 sky130_fd_sc_hd__a21o_1 _4122_ (.A1(_0755_),
    .A2(\tms1x00.A[1] ),
    .B1(_1992_),
    .X(_1994_));
 sky130_fd_sc_hd__o211a_1 _4123_ (.A1(net73),
    .A2(_1991_),
    .B1(_1994_),
    .C1(_1989_),
    .X(_0547_));
 sky130_fd_sc_hd__a21o_1 _4124_ (.A1(_0755_),
    .A2(\tms1x00.A[2] ),
    .B1(_1992_),
    .X(_1995_));
 sky130_fd_sc_hd__o211a_1 _4125_ (.A1(net74),
    .A2(_1991_),
    .B1(_1995_),
    .C1(_1989_),
    .X(_0548_));
 sky130_fd_sc_hd__a21o_1 _4126_ (.A1(_0755_),
    .A2(\tms1x00.A[3] ),
    .B1(_1992_),
    .X(_1996_));
 sky130_fd_sc_hd__o211a_1 _4127_ (.A1(net75),
    .A2(_1991_),
    .B1(_1996_),
    .C1(_1989_),
    .X(_0549_));
 sky130_fd_sc_hd__a21o_1 _4128_ (.A1(\tms1x00.status ),
    .A2(_0755_),
    .B1(_1992_),
    .X(_1997_));
 sky130_fd_sc_hd__o211a_1 _4129_ (.A1(net76),
    .A2(_1991_),
    .B1(_1997_),
    .C1(_1989_),
    .X(_0550_));
 sky130_fd_sc_hd__and3b_1 _4130_ (.A_N(net78),
    .B(net151),
    .C(net79),
    .X(_1998_));
 sky130_fd_sc_hd__nand2_2 _4131_ (.A(_1936_),
    .B(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__nand2_1 _4132_ (.A(\tms1x00.status ),
    .B(\tms1x00.ins_in[0] ),
    .Y(_2000_));
 sky130_fd_sc_hd__nor2_2 _4133_ (.A(_1999_),
    .B(_2000_),
    .Y(_2001_));
 sky130_fd_sc_hd__a21o_1 _4134_ (.A1(\tms1x00.ins_in[1] ),
    .A2(_2001_),
    .B1(\tms1x00.CL ),
    .X(_2002_));
 sky130_fd_sc_hd__or4_2 _4135_ (.A(_0748_),
    .B(_0744_),
    .C(_1135_),
    .D(_1999_),
    .X(_2003_));
 sky130_fd_sc_hd__and3_1 _4136_ (.A(_1922_),
    .B(_2002_),
    .C(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__clkbuf_1 _4137_ (.A(_2004_),
    .X(_0551_));
 sky130_fd_sc_hd__or3b_1 _4138_ (.A(\tms1x00.status ),
    .B(_1910_),
    .C_N(_1999_),
    .X(_2005_));
 sky130_fd_sc_hd__clkbuf_1 _4139_ (.A(_2005_),
    .X(_0552_));
 sky130_fd_sc_hd__and4b_1 _4140_ (.A_N(\tms1x00.CL ),
    .B(\tms1x00.ins_in[1] ),
    .C(_0718_),
    .D(_2001_),
    .X(_2006_));
 sky130_fd_sc_hd__buf_2 _4141_ (.A(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__mux2_1 _4142_ (.A0(\tms1x00.SR[0] ),
    .A1(\tms1x00.PC[0] ),
    .S(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__clkbuf_1 _4143_ (.A(_2008_),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _4144_ (.A0(\tms1x00.SR[1] ),
    .A1(\tms1x00.PC[1] ),
    .S(_2007_),
    .X(_2009_));
 sky130_fd_sc_hd__clkbuf_1 _4145_ (.A(_2009_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _4146_ (.A0(\tms1x00.SR[2] ),
    .A1(\tms1x00.PC[2] ),
    .S(_2007_),
    .X(_2010_));
 sky130_fd_sc_hd__clkbuf_1 _4147_ (.A(_2010_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _4148_ (.A0(\tms1x00.SR[3] ),
    .A1(\tms1x00.PC[3] ),
    .S(_2007_),
    .X(_2011_));
 sky130_fd_sc_hd__clkbuf_1 _4149_ (.A(_2011_),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _4150_ (.A0(\tms1x00.SR[4] ),
    .A1(\tms1x00.PC[4] ),
    .S(_2007_),
    .X(_2012_));
 sky130_fd_sc_hd__clkbuf_1 _4151_ (.A(_2012_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _4152_ (.A0(\tms1x00.SR[5] ),
    .A1(\tms1x00.PC[5] ),
    .S(_2007_),
    .X(_2013_));
 sky130_fd_sc_hd__clkbuf_1 _4153_ (.A(_2013_),
    .X(_0558_));
 sky130_fd_sc_hd__or3b_1 _4154_ (.A(_0910_),
    .B(\tms1x00.ins_in[2] ),
    .C_N(_0906_),
    .X(_2014_));
 sky130_fd_sc_hd__nor2_2 _4155_ (.A(_0746_),
    .B(_2014_),
    .Y(_2015_));
 sky130_fd_sc_hd__mux2_1 _4156_ (.A0(\tms1x00.PA[0] ),
    .A1(_0743_),
    .S(_2015_),
    .X(_2016_));
 sky130_fd_sc_hd__inv_2 _4157_ (.A(_2014_),
    .Y(_2017_));
 sky130_fd_sc_hd__a22o_2 _4158_ (.A1(\tms1x00.ins_in[1] ),
    .A2(_2001_),
    .B1(_2017_),
    .B2(_0757_),
    .X(_2018_));
 sky130_fd_sc_hd__mux2_1 _4159_ (.A0(\tms1x00.PB[0] ),
    .A1(_2016_),
    .S(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__or2_1 _4160_ (.A(_1910_),
    .B(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__clkbuf_1 _4161_ (.A(_2020_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _4162_ (.A0(\tms1x00.PA[1] ),
    .A1(_1928_),
    .S(_2015_),
    .X(_2021_));
 sky130_fd_sc_hd__mux2_1 _4163_ (.A0(\tms1x00.PB[1] ),
    .A1(_2021_),
    .S(_2018_),
    .X(_2022_));
 sky130_fd_sc_hd__or2_1 _4164_ (.A(_1910_),
    .B(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__clkbuf_1 _4165_ (.A(_2023_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _4166_ (.A0(\tms1x00.PA[2] ),
    .A1(\tms1x00.ins_in[6] ),
    .S(_2015_),
    .X(_2024_));
 sky130_fd_sc_hd__mux2_1 _4167_ (.A0(\tms1x00.PB[2] ),
    .A1(_2024_),
    .S(_2018_),
    .X(_2025_));
 sky130_fd_sc_hd__or2_1 _4168_ (.A(_1910_),
    .B(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__clkbuf_1 _4169_ (.A(_2026_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _4170_ (.A0(\tms1x00.PA[3] ),
    .A1(_0742_),
    .S(_2015_),
    .X(_2027_));
 sky130_fd_sc_hd__mux2_1 _4171_ (.A0(\tms1x00.PB[3] ),
    .A1(_2027_),
    .S(_2018_),
    .X(_2028_));
 sky130_fd_sc_hd__or2_1 _4172_ (.A(_1910_),
    .B(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__clkbuf_1 _4173_ (.A(_2029_),
    .X(_0562_));
 sky130_fd_sc_hd__o31ai_4 _4174_ (.A1(\tms1x00.CL ),
    .A2(_1999_),
    .A3(_2000_),
    .B1(_2003_),
    .Y(_2030_));
 sky130_fd_sc_hd__mux2_1 _4175_ (.A0(\tms1x00.PA[0] ),
    .A1(\tms1x00.PB[0] ),
    .S(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__or2_1 _4176_ (.A(_1910_),
    .B(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__clkbuf_1 _4177_ (.A(_2032_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _4178_ (.A0(\tms1x00.PA[1] ),
    .A1(\tms1x00.PB[1] ),
    .S(_2030_),
    .X(_2033_));
 sky130_fd_sc_hd__or2_1 _4179_ (.A(_1910_),
    .B(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__clkbuf_1 _4180_ (.A(_2034_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _4181_ (.A0(\tms1x00.PA[2] ),
    .A1(\tms1x00.PB[2] ),
    .S(_2030_),
    .X(_2035_));
 sky130_fd_sc_hd__or2_1 _4182_ (.A(_1910_),
    .B(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__clkbuf_1 _4183_ (.A(_2036_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _4184_ (.A0(\tms1x00.PA[3] ),
    .A1(\tms1x00.PB[3] ),
    .S(_2030_),
    .X(_2037_));
 sky130_fd_sc_hd__or2_1 _4185_ (.A(_1910_),
    .B(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__clkbuf_1 _4186_ (.A(_2038_),
    .X(_0566_));
 sky130_fd_sc_hd__or3_2 _4187_ (.A(net79),
    .B(net78),
    .C(_0723_),
    .X(_2039_));
 sky130_fd_sc_hd__nor2_2 _4188_ (.A(net151),
    .B(_2039_),
    .Y(_2040_));
 sky130_fd_sc_hd__nand2_1 _4189_ (.A(_0853_),
    .B(_0904_),
    .Y(_2041_));
 sky130_fd_sc_hd__and2_1 _4190_ (.A(_0911_),
    .B(_2017_),
    .X(_2042_));
 sky130_fd_sc_hd__nor2_1 _4191_ (.A(_2041_),
    .B(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__nand2_1 _4192_ (.A(\tms1x00.ins_in[1] ),
    .B(\tms1x00.ins_in[0] ),
    .Y(_2044_));
 sky130_fd_sc_hd__or2_1 _4193_ (.A(_0912_),
    .B(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__or4_1 _4194_ (.A(_0742_),
    .B(\tms1x00.ins_in[6] ),
    .C(_1928_),
    .D(_0743_),
    .X(_2046_));
 sky130_fd_sc_hd__nor2_1 _4195_ (.A(_0910_),
    .B(_2046_),
    .Y(_2047_));
 sky130_fd_sc_hd__a22o_1 _4196_ (.A1(_0743_),
    .A2(_1027_),
    .B1(_2047_),
    .B2(\tms1x00.K_latch[0] ),
    .X(_2048_));
 sky130_fd_sc_hd__or2_1 _4197_ (.A(net151),
    .B(_2039_),
    .X(_2049_));
 sky130_fd_sc_hd__a211o_1 _4198_ (.A1(\tms1x00.Y[0] ),
    .A2(_2045_),
    .B1(_2048_),
    .C1(_2049_),
    .X(_2050_));
 sky130_fd_sc_hd__o22a_1 _4199_ (.A1(\tms1x00.P[0] ),
    .A2(_2040_),
    .B1(_2043_),
    .B2(_2050_),
    .X(_0567_));
 sky130_fd_sc_hd__nand2_1 _4200_ (.A(_0980_),
    .B(_1026_),
    .Y(_2051_));
 sky130_fd_sc_hd__nor2_1 _4201_ (.A(_2051_),
    .B(_2042_),
    .Y(_2052_));
 sky130_fd_sc_hd__a22o_1 _4202_ (.A1(_1928_),
    .A2(_1027_),
    .B1(_2047_),
    .B2(\tms1x00.K_latch[1] ),
    .X(_2053_));
 sky130_fd_sc_hd__a211o_1 _4203_ (.A1(\tms1x00.Y[1] ),
    .A2(_2045_),
    .B1(_2053_),
    .C1(_2049_),
    .X(_2054_));
 sky130_fd_sc_hd__o22a_1 _4204_ (.A1(\tms1x00.P[1] ),
    .A2(_2040_),
    .B1(_2052_),
    .B2(_2054_),
    .X(_0568_));
 sky130_fd_sc_hd__nand2_1 _4205_ (.A(_1082_),
    .B(_1127_),
    .Y(_2055_));
 sky130_fd_sc_hd__nor2_1 _4206_ (.A(_2055_),
    .B(_2042_),
    .Y(_2056_));
 sky130_fd_sc_hd__a221o_1 _4207_ (.A1(\tms1x00.K_latch[2] ),
    .A2(_2047_),
    .B1(_2045_),
    .B2(_0729_),
    .C1(_1027_),
    .X(_2057_));
 sky130_fd_sc_hd__or2_1 _4208_ (.A(_2049_),
    .B(_2057_),
    .X(_2058_));
 sky130_fd_sc_hd__o22a_1 _4209_ (.A1(\tms1x00.P[2] ),
    .A2(_2040_),
    .B1(_2056_),
    .B2(_2058_),
    .X(_0569_));
 sky130_fd_sc_hd__nor2_1 _4210_ (.A(_1225_),
    .B(_2042_),
    .Y(_2059_));
 sky130_fd_sc_hd__a221o_1 _4211_ (.A1(\tms1x00.K_latch[3] ),
    .A2(_2047_),
    .B1(_2045_),
    .B2(_0732_),
    .C1(_2049_),
    .X(_2060_));
 sky130_fd_sc_hd__o22a_1 _4212_ (.A1(\tms1x00.P[3] ),
    .A2(_2040_),
    .B1(_2059_),
    .B2(_2060_),
    .X(_0570_));
 sky130_fd_sc_hd__and3_1 _4213_ (.A(\tms1x00.CL ),
    .B(_0758_),
    .C(_1136_),
    .X(_2061_));
 sky130_fd_sc_hd__a21o_1 _4214_ (.A1(\tms1x00.status ),
    .A2(\tms1x00.ins_in[0] ),
    .B1(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__nand2_1 _4215_ (.A(_1998_),
    .B(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__a32o_1 _4216_ (.A1(\tms1x00.status ),
    .A2(\tms1x00.ins_in[2] ),
    .A3(\tms1x00.ins_in[0] ),
    .B1(\tms1x00.SR[0] ),
    .B2(_2061_),
    .X(_2064_));
 sky130_fd_sc_hd__a22o_1 _4217_ (.A1(\tms1x00.PC[0] ),
    .A2(_2063_),
    .B1(_2064_),
    .B2(_1998_),
    .X(_2065_));
 sky130_fd_sc_hd__nor2_1 _4218_ (.A(\tms1x00.PC[0] ),
    .B(_0721_),
    .Y(_2066_));
 sky130_fd_sc_hd__a211o_1 _4219_ (.A1(_0721_),
    .A2(_2065_),
    .B1(_2066_),
    .C1(_0745_),
    .X(_2067_));
 sky130_fd_sc_hd__o211a_1 _4220_ (.A1(\tms1x00.PC[0] ),
    .A2(_1936_),
    .B1(_2067_),
    .C1(_1989_),
    .X(_0571_));
 sky130_fd_sc_hd__nand2_1 _4221_ (.A(\tms1x00.CL ),
    .B(\tms1x00.SR[1] ),
    .Y(_2068_));
 sky130_fd_sc_hd__o2bb2a_1 _4222_ (.A1_N(\tms1x00.ins_in[3] ),
    .A2_N(_2001_),
    .B1(_2003_),
    .B2(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__o21a_1 _4223_ (.A1(_0745_),
    .A2(_2063_),
    .B1(_1919_),
    .X(_2070_));
 sky130_fd_sc_hd__nand2_1 _4224_ (.A(\tms1x00.PC[1] ),
    .B(_2070_),
    .Y(_2071_));
 sky130_fd_sc_hd__a21oi_1 _4225_ (.A1(_2069_),
    .A2(_2071_),
    .B1(net106),
    .Y(_0572_));
 sky130_fd_sc_hd__and3_1 _4226_ (.A(_1936_),
    .B(_1998_),
    .C(_2061_),
    .X(_2072_));
 sky130_fd_sc_hd__a22o_1 _4227_ (.A1(_0743_),
    .A2(_2001_),
    .B1(_2072_),
    .B2(\tms1x00.SR[2] ),
    .X(_2073_));
 sky130_fd_sc_hd__a21oi_1 _4228_ (.A1(\tms1x00.PC[2] ),
    .A2(_2070_),
    .B1(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__nor2_1 _4229_ (.A(net106),
    .B(_2074_),
    .Y(_0573_));
 sky130_fd_sc_hd__a22o_1 _4230_ (.A1(_1928_),
    .A2(_2001_),
    .B1(_2072_),
    .B2(\tms1x00.SR[3] ),
    .X(_2075_));
 sky130_fd_sc_hd__a21oi_1 _4231_ (.A1(\tms1x00.PC[3] ),
    .A2(_2070_),
    .B1(_2075_),
    .Y(_2076_));
 sky130_fd_sc_hd__nor2_1 _4232_ (.A(net106),
    .B(_2076_),
    .Y(_0574_));
 sky130_fd_sc_hd__a22o_1 _4233_ (.A1(\tms1x00.ins_in[6] ),
    .A2(_2001_),
    .B1(_2072_),
    .B2(\tms1x00.SR[4] ),
    .X(_2077_));
 sky130_fd_sc_hd__a21oi_1 _4234_ (.A1(\tms1x00.PC[4] ),
    .A2(_2070_),
    .B1(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hd__nor2_1 _4235_ (.A(net106),
    .B(_2078_),
    .Y(_0575_));
 sky130_fd_sc_hd__a22o_1 _4236_ (.A1(_0742_),
    .A2(_2001_),
    .B1(_2072_),
    .B2(\tms1x00.SR[5] ),
    .X(_2079_));
 sky130_fd_sc_hd__a21oi_1 _4237_ (.A1(\tms1x00.PC[5] ),
    .A2(_2070_),
    .B1(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__nor2_1 _4238_ (.A(net106),
    .B(_2080_),
    .Y(_0576_));
 sky130_fd_sc_hd__or2b_1 _4239_ (.A(\tms1x00.ins_in[6] ),
    .B_N(_0742_),
    .X(_2081_));
 sky130_fd_sc_hd__or4_1 _4240_ (.A(\tms1x00.ins_in[5] ),
    .B(_0743_),
    .C(\tms1x00.N[0] ),
    .D(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__o31ai_1 _4241_ (.A1(_1928_),
    .A2(_0743_),
    .A3(_2081_),
    .B1(\tms1x00.N[0] ),
    .Y(_2083_));
 sky130_fd_sc_hd__and2_1 _4242_ (.A(_2082_),
    .B(_2083_),
    .X(_2084_));
 sky130_fd_sc_hd__xor2_1 _4243_ (.A(\tms1x00.P[0] ),
    .B(_2084_),
    .X(_2085_));
 sky130_fd_sc_hd__and3_1 _4244_ (.A(_1928_),
    .B(_0756_),
    .C(_0925_),
    .X(_2086_));
 sky130_fd_sc_hd__clkbuf_2 _4245_ (.A(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__mux2_1 _4246_ (.A0(\tms1x00.Y[0] ),
    .A1(_2085_),
    .S(_2087_),
    .X(_2088_));
 sky130_fd_sc_hd__and2_1 _4247_ (.A(_0762_),
    .B(_2088_),
    .X(_2089_));
 sky130_fd_sc_hd__clkbuf_1 _4248_ (.A(_2089_),
    .X(_0577_));
 sky130_fd_sc_hd__and2_1 _4249_ (.A(\tms1x00.P[1] ),
    .B(\tms1x00.N[1] ),
    .X(_2090_));
 sky130_fd_sc_hd__nor2_1 _4250_ (.A(\tms1x00.P[1] ),
    .B(\tms1x00.N[1] ),
    .Y(_2091_));
 sky130_fd_sc_hd__or2_1 _4251_ (.A(_2090_),
    .B(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__a21boi_1 _4252_ (.A1(\tms1x00.P[0] ),
    .A2(_2082_),
    .B1_N(_2083_),
    .Y(_2093_));
 sky130_fd_sc_hd__xnor2_1 _4253_ (.A(_2092_),
    .B(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__nand2_1 _4254_ (.A(_2087_),
    .B(_2094_),
    .Y(_2095_));
 sky130_fd_sc_hd__o211a_1 _4255_ (.A1(\tms1x00.Y[1] ),
    .A2(_2087_),
    .B1(_2095_),
    .C1(_1989_),
    .X(_0578_));
 sky130_fd_sc_hd__nand2_1 _4256_ (.A(\tms1x00.P[2] ),
    .B(\tms1x00.N[2] ),
    .Y(_2096_));
 sky130_fd_sc_hd__or2_1 _4257_ (.A(\tms1x00.P[2] ),
    .B(\tms1x00.N[2] ),
    .X(_2097_));
 sky130_fd_sc_hd__nand2_1 _4258_ (.A(_2096_),
    .B(_2097_),
    .Y(_2098_));
 sky130_fd_sc_hd__o21ba_1 _4259_ (.A1(_2091_),
    .A2(_2093_),
    .B1_N(_2090_),
    .X(_2099_));
 sky130_fd_sc_hd__xnor2_1 _4260_ (.A(_2098_),
    .B(_2099_),
    .Y(_2100_));
 sky130_fd_sc_hd__nand2_1 _4261_ (.A(_2087_),
    .B(_2100_),
    .Y(_2101_));
 sky130_fd_sc_hd__o211a_1 _4262_ (.A1(_0729_),
    .A2(_2087_),
    .B1(_2101_),
    .C1(_1989_),
    .X(_0579_));
 sky130_fd_sc_hd__o21ai_1 _4263_ (.A1(_2098_),
    .A2(_2099_),
    .B1(_2096_),
    .Y(_2102_));
 sky130_fd_sc_hd__xor2_1 _4264_ (.A(\tms1x00.P[3] ),
    .B(\tms1x00.N[3] ),
    .X(_2103_));
 sky130_fd_sc_hd__xnor2_1 _4265_ (.A(_2102_),
    .B(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__nand2_1 _4266_ (.A(_2087_),
    .B(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__o211a_1 _4267_ (.A1(_0733_),
    .A2(_2087_),
    .B1(_2105_),
    .C1(_1989_),
    .X(_0580_));
 sky130_fd_sc_hd__and3_1 _4268_ (.A(_1928_),
    .B(_0743_),
    .C(_0907_),
    .X(_2106_));
 sky130_fd_sc_hd__nor2_1 _4269_ (.A(_0748_),
    .B(_2046_),
    .Y(_2107_));
 sky130_fd_sc_hd__o21a_1 _4270_ (.A1(_2106_),
    .A2(_2107_),
    .B1(_0757_),
    .X(_2108_));
 sky130_fd_sc_hd__mux2_1 _4271_ (.A0(\tms1x00.X[0] ),
    .A1(_0763_),
    .S(_2106_),
    .X(_2109_));
 sky130_fd_sc_hd__nand2_1 _4272_ (.A(_2108_),
    .B(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__o211a_1 _4273_ (.A1(\tms1x00.X[0] ),
    .A2(_2108_),
    .B1(_2110_),
    .C1(_0762_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _4274_ (.A0(\tms1x00.X[1] ),
    .A1(_0755_),
    .S(_2106_),
    .X(_2111_));
 sky130_fd_sc_hd__nand2_1 _4275_ (.A(_2108_),
    .B(_2111_),
    .Y(_2112_));
 sky130_fd_sc_hd__o211a_1 _4276_ (.A1(\tms1x00.X[1] ),
    .A2(_2108_),
    .B1(_2112_),
    .C1(_0762_),
    .X(_0582_));
 sky130_fd_sc_hd__o21ai_1 _4277_ (.A1(\tms1x00.X[2] ),
    .A2(_1928_),
    .B1(_2108_),
    .Y(_2113_));
 sky130_fd_sc_hd__o211a_1 _4278_ (.A1(\tms1x00.X[2] ),
    .A2(_2108_),
    .B1(_2113_),
    .C1(_0762_),
    .X(_0583_));
 sky130_fd_sc_hd__or2_1 _4279_ (.A(\tms1x00.N[0] ),
    .B(_2040_),
    .X(_2114_));
 sky130_fd_sc_hd__clkbuf_1 _4280_ (.A(_2114_),
    .X(_0584_));
 sky130_fd_sc_hd__or2_1 _4281_ (.A(\tms1x00.N[1] ),
    .B(_2040_),
    .X(_2115_));
 sky130_fd_sc_hd__clkbuf_1 _4282_ (.A(_2115_),
    .X(_0585_));
 sky130_fd_sc_hd__or2_1 _4283_ (.A(\tms1x00.N[2] ),
    .B(_2040_),
    .X(_2116_));
 sky130_fd_sc_hd__clkbuf_1 _4284_ (.A(_2116_),
    .X(_0586_));
 sky130_fd_sc_hd__or2_1 _4285_ (.A(\tms1x00.N[3] ),
    .B(_2040_),
    .X(_2117_));
 sky130_fd_sc_hd__clkbuf_1 _4286_ (.A(_2117_),
    .X(_0587_));
 sky130_fd_sc_hd__or4b_1 _4287_ (.A(_0723_),
    .B(_2081_),
    .C(_0746_),
    .D_N(_1990_),
    .X(_2118_));
 sky130_fd_sc_hd__clkbuf_2 _4288_ (.A(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__mux2_1 _4289_ (.A0(_2085_),
    .A1(\tms1x00.A[0] ),
    .S(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__clkbuf_1 _4290_ (.A(_2120_),
    .X(_0588_));
 sky130_fd_sc_hd__nand2_1 _4291_ (.A(\tms1x00.A[1] ),
    .B(_2119_),
    .Y(_2121_));
 sky130_fd_sc_hd__o21ai_1 _4292_ (.A1(_2094_),
    .A2(_2119_),
    .B1(_2121_),
    .Y(_0589_));
 sky130_fd_sc_hd__nand2_1 _4293_ (.A(\tms1x00.A[2] ),
    .B(_2119_),
    .Y(_2122_));
 sky130_fd_sc_hd__o21ai_1 _4294_ (.A1(_2100_),
    .A2(_2119_),
    .B1(_2122_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _4295_ (.A(\tms1x00.A[3] ),
    .B(_2119_),
    .Y(_2123_));
 sky130_fd_sc_hd__o21ai_1 _4296_ (.A1(_2104_),
    .A2(_2119_),
    .B1(_2123_),
    .Y(_0591_));
 sky130_fd_sc_hd__nor2_2 _4297_ (.A(_1316_),
    .B(_1397_),
    .Y(_2124_));
 sky130_fd_sc_hd__mux2_1 _4298_ (.A0(\tms1x00.RAM[119][0] ),
    .A1(_1335_),
    .S(_2124_),
    .X(_2125_));
 sky130_fd_sc_hd__clkbuf_1 _4299_ (.A(_2125_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(\tms1x00.RAM[119][1] ),
    .A1(_1342_),
    .S(_2124_),
    .X(_2126_));
 sky130_fd_sc_hd__clkbuf_1 _4301_ (.A(_2126_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(\tms1x00.RAM[119][2] ),
    .A1(_1345_),
    .S(_2124_),
    .X(_2127_));
 sky130_fd_sc_hd__clkbuf_1 _4303_ (.A(_2127_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _4304_ (.A0(\tms1x00.RAM[119][3] ),
    .A1(_1348_),
    .S(_2124_),
    .X(_2128_));
 sky130_fd_sc_hd__clkbuf_1 _4305_ (.A(_2128_),
    .X(_0595_));
 sky130_fd_sc_hd__nor2_2 _4306_ (.A(_1697_),
    .B(_1534_),
    .Y(_2129_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(\tms1x00.RAM[39][0] ),
    .A1(_1335_),
    .S(_2129_),
    .X(_2130_));
 sky130_fd_sc_hd__clkbuf_1 _4308_ (.A(_2130_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(\tms1x00.RAM[39][1] ),
    .A1(_1342_),
    .S(_2129_),
    .X(_2131_));
 sky130_fd_sc_hd__clkbuf_1 _4310_ (.A(_2131_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(\tms1x00.RAM[39][2] ),
    .A1(_1345_),
    .S(_2129_),
    .X(_2132_));
 sky130_fd_sc_hd__clkbuf_1 _4312_ (.A(_2132_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(\tms1x00.RAM[39][3] ),
    .A1(_1348_),
    .S(_2129_),
    .X(_2133_));
 sky130_fd_sc_hd__clkbuf_1 _4314_ (.A(_2133_),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_2 _4315_ (.A(_1241_),
    .B(_1324_),
    .Y(_2134_));
 sky130_fd_sc_hd__mux2_1 _4316_ (.A0(\tms1x00.RAM[22][0] ),
    .A1(_1335_),
    .S(_2134_),
    .X(_2135_));
 sky130_fd_sc_hd__clkbuf_1 _4317_ (.A(_2135_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _4318_ (.A0(\tms1x00.RAM[22][1] ),
    .A1(_1342_),
    .S(_2134_),
    .X(_2136_));
 sky130_fd_sc_hd__clkbuf_1 _4319_ (.A(_2136_),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(\tms1x00.RAM[22][2] ),
    .A1(_1345_),
    .S(_2134_),
    .X(_2137_));
 sky130_fd_sc_hd__clkbuf_1 _4321_ (.A(_2137_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _4322_ (.A0(\tms1x00.RAM[22][3] ),
    .A1(_1348_),
    .S(_2134_),
    .X(_2138_));
 sky130_fd_sc_hd__clkbuf_1 _4323_ (.A(_2138_),
    .X(_0603_));
 sky130_fd_sc_hd__nor2_2 _4324_ (.A(_0928_),
    .B(_1241_),
    .Y(_2139_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(\tms1x00.RAM[29][0] ),
    .A1(_1335_),
    .S(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__clkbuf_1 _4326_ (.A(_2140_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _4327_ (.A0(\tms1x00.RAM[29][1] ),
    .A1(_1342_),
    .S(_2139_),
    .X(_2141_));
 sky130_fd_sc_hd__clkbuf_1 _4328_ (.A(_2141_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _4329_ (.A0(\tms1x00.RAM[29][2] ),
    .A1(_1345_),
    .S(_2139_),
    .X(_2142_));
 sky130_fd_sc_hd__clkbuf_1 _4330_ (.A(_2142_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(\tms1x00.RAM[29][3] ),
    .A1(_1348_),
    .S(_2139_),
    .X(_2143_));
 sky130_fd_sc_hd__clkbuf_1 _4332_ (.A(_2143_),
    .X(_0607_));
 sky130_fd_sc_hd__or2_2 _4333_ (.A(_1240_),
    .B(_1278_),
    .X(_2144_));
 sky130_fd_sc_hd__mux2_1 _4334_ (.A0(_1867_),
    .A1(\tms1x00.RAM[21][0] ),
    .S(_2144_),
    .X(_2145_));
 sky130_fd_sc_hd__clkbuf_1 _4335_ (.A(_2145_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(_1870_),
    .A1(\tms1x00.RAM[21][1] ),
    .S(_2144_),
    .X(_2146_));
 sky130_fd_sc_hd__clkbuf_1 _4337_ (.A(_2146_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(_1872_),
    .A1(\tms1x00.RAM[21][2] ),
    .S(_2144_),
    .X(_2147_));
 sky130_fd_sc_hd__clkbuf_1 _4339_ (.A(_2147_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _4340_ (.A0(_1874_),
    .A1(\tms1x00.RAM[21][3] ),
    .S(_2144_),
    .X(_2148_));
 sky130_fd_sc_hd__clkbuf_1 _4341_ (.A(_2148_),
    .X(_0611_));
 sky130_fd_sc_hd__or2_1 _4342_ (.A(_1242_),
    .B(_1240_),
    .X(_2149_));
 sky130_fd_sc_hd__or2_2 _4343_ (.A(_2149_),
    .B(_1353_),
    .X(_2150_));
 sky130_fd_sc_hd__mux2_1 _4344_ (.A0(_1867_),
    .A1(\tms1x00.RAM[16][0] ),
    .S(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__clkbuf_1 _4345_ (.A(_2151_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _4346_ (.A0(_1870_),
    .A1(\tms1x00.RAM[16][1] ),
    .S(_2150_),
    .X(_2152_));
 sky130_fd_sc_hd__clkbuf_1 _4347_ (.A(_2152_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _4348_ (.A0(_1872_),
    .A1(\tms1x00.RAM[16][2] ),
    .S(_2150_),
    .X(_2153_));
 sky130_fd_sc_hd__clkbuf_1 _4349_ (.A(_2153_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _4350_ (.A0(_1874_),
    .A1(\tms1x00.RAM[16][3] ),
    .S(_2150_),
    .X(_2154_));
 sky130_fd_sc_hd__clkbuf_1 _4351_ (.A(_2154_),
    .X(_0615_));
 sky130_fd_sc_hd__or2_4 _4352_ (.A(_2149_),
    .B(_1337_),
    .X(_2155_));
 sky130_fd_sc_hd__mux2_1 _4353_ (.A0(_1867_),
    .A1(\tms1x00.RAM[20][0] ),
    .S(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__clkbuf_1 _4354_ (.A(_2156_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _4355_ (.A0(_1870_),
    .A1(\tms1x00.RAM[20][1] ),
    .S(_2155_),
    .X(_2157_));
 sky130_fd_sc_hd__clkbuf_1 _4356_ (.A(_2157_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _4357_ (.A0(_1872_),
    .A1(\tms1x00.RAM[20][2] ),
    .S(_2155_),
    .X(_2158_));
 sky130_fd_sc_hd__clkbuf_1 _4358_ (.A(_2158_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _4359_ (.A0(_1874_),
    .A1(\tms1x00.RAM[20][3] ),
    .S(_2155_),
    .X(_2159_));
 sky130_fd_sc_hd__clkbuf_1 _4360_ (.A(_2159_),
    .X(_0619_));
 sky130_fd_sc_hd__or2_2 _4361_ (.A(_1352_),
    .B(_1422_),
    .X(_2160_));
 sky130_fd_sc_hd__mux2_1 _4362_ (.A0(_1867_),
    .A1(\tms1x00.RAM[12][0] ),
    .S(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__clkbuf_1 _4363_ (.A(_2161_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _4364_ (.A0(_1870_),
    .A1(\tms1x00.RAM[12][1] ),
    .S(_2160_),
    .X(_2162_));
 sky130_fd_sc_hd__clkbuf_1 _4365_ (.A(_2162_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _4366_ (.A0(_1872_),
    .A1(\tms1x00.RAM[12][2] ),
    .S(_2160_),
    .X(_2163_));
 sky130_fd_sc_hd__clkbuf_1 _4367_ (.A(_2163_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _4368_ (.A0(_1874_),
    .A1(\tms1x00.RAM[12][3] ),
    .S(_2160_),
    .X(_2164_));
 sky130_fd_sc_hd__clkbuf_1 _4369_ (.A(_2164_),
    .X(_0623_));
 sky130_fd_sc_hd__or2_2 _4370_ (.A(_1261_),
    .B(_1397_),
    .X(_2165_));
 sky130_fd_sc_hd__mux2_1 _4371_ (.A0(_1867_),
    .A1(\tms1x00.RAM[127][0] ),
    .S(_2165_),
    .X(_2166_));
 sky130_fd_sc_hd__clkbuf_1 _4372_ (.A(_2166_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _4373_ (.A0(_1870_),
    .A1(\tms1x00.RAM[127][1] ),
    .S(_2165_),
    .X(_2167_));
 sky130_fd_sc_hd__clkbuf_1 _4374_ (.A(_2167_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _4375_ (.A0(_1872_),
    .A1(\tms1x00.RAM[127][2] ),
    .S(_2165_),
    .X(_2168_));
 sky130_fd_sc_hd__clkbuf_1 _4376_ (.A(_2168_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _4377_ (.A0(_1874_),
    .A1(\tms1x00.RAM[127][3] ),
    .S(_2165_),
    .X(_2169_));
 sky130_fd_sc_hd__clkbuf_1 _4378_ (.A(_2169_),
    .X(_0627_));
 sky130_fd_sc_hd__or2_2 _4379_ (.A(_1261_),
    .B(_1473_),
    .X(_2170_));
 sky130_fd_sc_hd__mux2_1 _4380_ (.A0(_0920_),
    .A1(\tms1x00.RAM[15][0] ),
    .S(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__clkbuf_1 _4381_ (.A(_2171_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _4382_ (.A0(_1032_),
    .A1(\tms1x00.RAM[15][1] ),
    .S(_2170_),
    .X(_2172_));
 sky130_fd_sc_hd__clkbuf_1 _4383_ (.A(_2172_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _4384_ (.A0(_1133_),
    .A1(\tms1x00.RAM[15][2] ),
    .S(_2170_),
    .X(_2173_));
 sky130_fd_sc_hd__clkbuf_1 _4385_ (.A(_2173_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _4386_ (.A0(_1229_),
    .A1(\tms1x00.RAM[15][3] ),
    .S(_2170_),
    .X(_2174_));
 sky130_fd_sc_hd__clkbuf_1 _4387_ (.A(_2174_),
    .X(_0631_));
 sky130_fd_sc_hd__or2_2 _4388_ (.A(_1243_),
    .B(_1352_),
    .X(_2175_));
 sky130_fd_sc_hd__mux2_1 _4389_ (.A0(_0920_),
    .A1(\tms1x00.RAM[1][0] ),
    .S(_2175_),
    .X(_2176_));
 sky130_fd_sc_hd__clkbuf_1 _4390_ (.A(_2176_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _4391_ (.A0(_1032_),
    .A1(\tms1x00.RAM[1][1] ),
    .S(_2175_),
    .X(_2177_));
 sky130_fd_sc_hd__clkbuf_1 _4392_ (.A(_2177_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _4393_ (.A0(_1133_),
    .A1(\tms1x00.RAM[1][2] ),
    .S(_2175_),
    .X(_2178_));
 sky130_fd_sc_hd__clkbuf_1 _4394_ (.A(_2178_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _4395_ (.A0(_1229_),
    .A1(\tms1x00.RAM[1][3] ),
    .S(_2175_),
    .X(_2179_));
 sky130_fd_sc_hd__clkbuf_1 _4396_ (.A(_2179_),
    .X(_0635_));
 sky130_fd_sc_hd__nor2_2 _4397_ (.A(_0928_),
    .B(_1352_),
    .Y(_2180_));
 sky130_fd_sc_hd__mux2_1 _4398_ (.A0(\tms1x00.RAM[13][0] ),
    .A1(_1335_),
    .S(_2180_),
    .X(_2181_));
 sky130_fd_sc_hd__clkbuf_1 _4399_ (.A(_2181_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _4400_ (.A0(\tms1x00.RAM[13][1] ),
    .A1(_1342_),
    .S(_2180_),
    .X(_2182_));
 sky130_fd_sc_hd__clkbuf_1 _4401_ (.A(_2182_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _4402_ (.A0(\tms1x00.RAM[13][2] ),
    .A1(_1345_),
    .S(_2180_),
    .X(_2183_));
 sky130_fd_sc_hd__clkbuf_1 _4403_ (.A(_2183_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _4404_ (.A0(\tms1x00.RAM[13][3] ),
    .A1(_1348_),
    .S(_2180_),
    .X(_2184_));
 sky130_fd_sc_hd__clkbuf_1 _4405_ (.A(_2184_),
    .X(_0639_));
 sky130_fd_sc_hd__or2_2 _4406_ (.A(_1352_),
    .B(_1410_),
    .X(_2185_));
 sky130_fd_sc_hd__mux2_1 _4407_ (.A0(_0920_),
    .A1(\tms1x00.RAM[14][0] ),
    .S(_2185_),
    .X(_2186_));
 sky130_fd_sc_hd__clkbuf_1 _4408_ (.A(_2186_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _4409_ (.A0(_1032_),
    .A1(\tms1x00.RAM[14][1] ),
    .S(_2185_),
    .X(_2187_));
 sky130_fd_sc_hd__clkbuf_1 _4410_ (.A(_2187_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _4411_ (.A0(_1133_),
    .A1(\tms1x00.RAM[14][2] ),
    .S(_2185_),
    .X(_2188_));
 sky130_fd_sc_hd__clkbuf_1 _4412_ (.A(_2188_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _4413_ (.A0(_1229_),
    .A1(\tms1x00.RAM[14][3] ),
    .S(_2185_),
    .X(_2189_));
 sky130_fd_sc_hd__clkbuf_1 _4414_ (.A(_2189_),
    .X(_0643_));
 sky130_fd_sc_hd__or2_2 _4415_ (.A(_1255_),
    .B(_1352_),
    .X(_2190_));
 sky130_fd_sc_hd__mux2_1 _4416_ (.A0(_0920_),
    .A1(\tms1x00.RAM[9][0] ),
    .S(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__clkbuf_1 _4417_ (.A(_2191_),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _4418_ (.A0(_1032_),
    .A1(\tms1x00.RAM[9][1] ),
    .S(_2190_),
    .X(_2192_));
 sky130_fd_sc_hd__clkbuf_1 _4419_ (.A(_2192_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _4420_ (.A0(_1133_),
    .A1(\tms1x00.RAM[9][2] ),
    .S(_2190_),
    .X(_2193_));
 sky130_fd_sc_hd__clkbuf_1 _4421_ (.A(_2193_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _4422_ (.A0(_1229_),
    .A1(\tms1x00.RAM[9][3] ),
    .S(_2190_),
    .X(_2194_));
 sky130_fd_sc_hd__clkbuf_1 _4423_ (.A(_2194_),
    .X(_0647_));
 sky130_fd_sc_hd__clkbuf_4 _4424_ (.A(_2039_),
    .X(_2195_));
 sky130_fd_sc_hd__mux2_1 _4425_ (.A0(\tms1x00.PC[0] ),
    .A1(\tms1x00.rom_addr[0] ),
    .S(_2195_),
    .X(_2196_));
 sky130_fd_sc_hd__clkbuf_1 _4426_ (.A(_2196_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _4427_ (.A0(\tms1x00.PC[1] ),
    .A1(\tms1x00.rom_addr[1] ),
    .S(_2195_),
    .X(_2197_));
 sky130_fd_sc_hd__clkbuf_1 _4428_ (.A(_2197_),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _4429_ (.A0(\tms1x00.PC[2] ),
    .A1(net98),
    .S(_2195_),
    .X(_2198_));
 sky130_fd_sc_hd__clkbuf_1 _4430_ (.A(_2198_),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _4431_ (.A0(\tms1x00.PC[3] ),
    .A1(net99),
    .S(_2195_),
    .X(_2199_));
 sky130_fd_sc_hd__clkbuf_1 _4432_ (.A(_2199_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _4433_ (.A0(\tms1x00.PC[4] ),
    .A1(net100),
    .S(_2195_),
    .X(_2200_));
 sky130_fd_sc_hd__clkbuf_1 _4434_ (.A(_2200_),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _4435_ (.A0(\tms1x00.PC[5] ),
    .A1(net101),
    .S(_2195_),
    .X(_2201_));
 sky130_fd_sc_hd__clkbuf_1 _4436_ (.A(_2201_),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _4437_ (.A0(\tms1x00.PA[0] ),
    .A1(net102),
    .S(_2195_),
    .X(_2202_));
 sky130_fd_sc_hd__clkbuf_1 _4438_ (.A(_2202_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _4439_ (.A0(\tms1x00.PA[1] ),
    .A1(net103),
    .S(_2195_),
    .X(_2203_));
 sky130_fd_sc_hd__clkbuf_1 _4440_ (.A(_2203_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _4441_ (.A0(\tms1x00.PA[2] ),
    .A1(net104),
    .S(_2195_),
    .X(_2204_));
 sky130_fd_sc_hd__clkbuf_1 _4442_ (.A(_2204_),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _4443_ (.A0(\tms1x00.PA[3] ),
    .A1(net105),
    .S(_2195_),
    .X(_2205_));
 sky130_fd_sc_hd__clkbuf_1 _4444_ (.A(_2205_),
    .X(_0657_));
 sky130_fd_sc_hd__dfxtp_2 _4445_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0049_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_4 _4446_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0000_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_2 _4447_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0002_),
    .Q(\tms1x00.wb_step ));
 sky130_fd_sc_hd__dfxtp_1 _4448_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0001_),
    .Q(wb_rst_override));
 sky130_fd_sc_hd__dfxtp_1 _4449_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0050_),
    .Q(chip_sel_override));
 sky130_fd_sc_hd__dfxtp_1 _4450_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0003_),
    .Q(\wbs_o_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4451_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0014_),
    .Q(\wbs_o_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4452_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0025_),
    .Q(\wbs_o_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4453_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0028_),
    .Q(\wbs_o_buff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4454_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0029_),
    .Q(\wbs_o_buff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4455_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0030_),
    .Q(\wbs_o_buff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4456_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0031_),
    .Q(\wbs_o_buff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4457_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0032_),
    .Q(\wbs_o_buff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4458_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0033_),
    .Q(\wbs_o_buff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4459_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0034_),
    .Q(\wbs_o_buff[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4460_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0004_),
    .Q(\wbs_o_buff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4461_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0005_),
    .Q(\wbs_o_buff[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4462_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0006_),
    .Q(\wbs_o_buff[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4463_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0007_),
    .Q(\wbs_o_buff[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4464_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0008_),
    .Q(\wbs_o_buff[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4465_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0009_),
    .Q(\wbs_o_buff[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4466_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0010_),
    .Q(\wbs_o_buff[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4467_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0011_),
    .Q(\wbs_o_buff[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4468_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0012_),
    .Q(\wbs_o_buff[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4469_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0013_),
    .Q(\wbs_o_buff[19] ));
 sky130_fd_sc_hd__dfxtp_1 _4470_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0015_),
    .Q(\wbs_o_buff[20] ));
 sky130_fd_sc_hd__dfxtp_1 _4471_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0016_),
    .Q(\wbs_o_buff[21] ));
 sky130_fd_sc_hd__dfxtp_1 _4472_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0017_),
    .Q(\wbs_o_buff[22] ));
 sky130_fd_sc_hd__dfxtp_1 _4473_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0018_),
    .Q(\wbs_o_buff[23] ));
 sky130_fd_sc_hd__dfxtp_1 _4474_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0019_),
    .Q(\wbs_o_buff[24] ));
 sky130_fd_sc_hd__dfxtp_1 _4475_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0020_),
    .Q(\wbs_o_buff[25] ));
 sky130_fd_sc_hd__dfxtp_1 _4476_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0021_),
    .Q(\wbs_o_buff[26] ));
 sky130_fd_sc_hd__dfxtp_1 _4477_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0022_),
    .Q(\wbs_o_buff[27] ));
 sky130_fd_sc_hd__dfxtp_1 _4478_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0023_),
    .Q(\wbs_o_buff[28] ));
 sky130_fd_sc_hd__dfxtp_1 _4479_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0024_),
    .Q(\wbs_o_buff[29] ));
 sky130_fd_sc_hd__dfxtp_1 _4480_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0026_),
    .Q(\wbs_o_buff[30] ));
 sky130_fd_sc_hd__dfxtp_1 _4481_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0027_),
    .Q(\wbs_o_buff[31] ));
 sky130_fd_sc_hd__dfxtp_1 _4482_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net204),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_1 _4483_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(valid),
    .Q(feedback_delay));
 sky130_fd_sc_hd__dfxtp_1 _4484_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0051_),
    .Q(\tms1x00.RAM[109][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4485_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0052_),
    .Q(\tms1x00.RAM[109][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4486_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0053_),
    .Q(\tms1x00.RAM[109][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4487_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0054_),
    .Q(\tms1x00.RAM[109][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4488_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0055_),
    .Q(\tms1x00.RAM[99][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4489_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0056_),
    .Q(\tms1x00.RAM[99][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4490_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0057_),
    .Q(\tms1x00.RAM[99][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4491_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0058_),
    .Q(\tms1x00.RAM[99][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4492_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0059_),
    .Q(\tms1x00.RAM[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4493_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0060_),
    .Q(\tms1x00.RAM[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4494_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0061_),
    .Q(\tms1x00.RAM[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4495_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0062_),
    .Q(\tms1x00.RAM[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4496_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0063_),
    .Q(\tms1x00.RAM[89][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4497_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0064_),
    .Q(\tms1x00.RAM[89][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4498_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0065_),
    .Q(\tms1x00.RAM[89][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4499_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0066_),
    .Q(\tms1x00.RAM[89][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4500_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0067_),
    .Q(\tms1x00.RAM[79][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4501_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0068_),
    .Q(\tms1x00.RAM[79][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4502_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0069_),
    .Q(\tms1x00.RAM[79][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4503_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0070_),
    .Q(\tms1x00.RAM[79][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4504_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0071_),
    .Q(\tms1x00.RAM[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4505_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0072_),
    .Q(\tms1x00.RAM[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4506_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0073_),
    .Q(\tms1x00.RAM[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4507_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0074_),
    .Q(\tms1x00.RAM[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4508_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0075_),
    .Q(\tms1x00.RAM[69][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4509_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0076_),
    .Q(\tms1x00.RAM[69][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4510_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0077_),
    .Q(\tms1x00.RAM[69][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4511_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0078_),
    .Q(\tms1x00.RAM[69][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4512_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0079_),
    .Q(\tms1x00.RAM[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4513_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0080_),
    .Q(\tms1x00.RAM[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4514_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0081_),
    .Q(\tms1x00.RAM[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4515_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0082_),
    .Q(\tms1x00.RAM[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4516_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0083_),
    .Q(\K_override[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4517_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0084_),
    .Q(\K_override[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4518_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0085_),
    .Q(\K_override[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4519_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0086_),
    .Q(\K_override[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4520_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0087_),
    .Q(\tms1x00.RAM[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4521_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0088_),
    .Q(\tms1x00.RAM[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4522_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0089_),
    .Q(\tms1x00.RAM[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4523_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0090_),
    .Q(\tms1x00.RAM[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4524_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0091_),
    .Q(\tms1x00.RAM[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4525_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0092_),
    .Q(\tms1x00.RAM[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4526_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0093_),
    .Q(\tms1x00.RAM[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4527_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0094_),
    .Q(\tms1x00.RAM[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4528_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0095_),
    .Q(\tms1x00.RAM[104][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4529_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0096_),
    .Q(\tms1x00.RAM[104][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4530_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0097_),
    .Q(\tms1x00.RAM[104][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4531_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0098_),
    .Q(\tms1x00.RAM[104][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4532_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0099_),
    .Q(\tms1x00.RAM[103][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4533_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0100_),
    .Q(\tms1x00.RAM[103][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4534_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0101_),
    .Q(\tms1x00.RAM[103][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4535_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0102_),
    .Q(\tms1x00.RAM[103][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4536_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0103_),
    .Q(\tms1x00.RAM[102][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4537_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0104_),
    .Q(\tms1x00.RAM[102][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4538_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0105_),
    .Q(\tms1x00.RAM[102][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4539_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0106_),
    .Q(\tms1x00.RAM[102][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4540_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0107_),
    .Q(\tms1x00.RAM[101][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4541_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0108_),
    .Q(\tms1x00.RAM[101][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4542_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0109_),
    .Q(\tms1x00.RAM[101][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4543_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0110_),
    .Q(\tms1x00.RAM[101][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4544_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0111_),
    .Q(\tms1x00.RAM[100][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4545_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0112_),
    .Q(\tms1x00.RAM[100][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4546_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0113_),
    .Q(\tms1x00.RAM[100][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4547_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0114_),
    .Q(\tms1x00.RAM[100][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4548_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0115_),
    .Q(\tms1x00.RAM[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4549_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0116_),
    .Q(\tms1x00.RAM[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4550_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0117_),
    .Q(\tms1x00.RAM[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4551_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0118_),
    .Q(\tms1x00.RAM[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4552_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0119_),
    .Q(\tms1x00.RAM[98][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4553_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0120_),
    .Q(\tms1x00.RAM[98][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4554_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0121_),
    .Q(\tms1x00.RAM[98][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4555_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0122_),
    .Q(\tms1x00.RAM[98][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4556_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0123_),
    .Q(\tms1x00.RAM[97][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4557_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0124_),
    .Q(\tms1x00.RAM[97][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4558_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0125_),
    .Q(\tms1x00.RAM[97][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4559_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0126_),
    .Q(\tms1x00.RAM[97][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4560_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0127_),
    .Q(\tms1x00.RAM[96][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4561_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0128_),
    .Q(\tms1x00.RAM[96][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4562_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0129_),
    .Q(\tms1x00.RAM[96][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4563_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0130_),
    .Q(\tms1x00.RAM[96][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4564_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0131_),
    .Q(\tms1x00.RAM[95][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4565_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0132_),
    .Q(\tms1x00.RAM[95][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4566_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0133_),
    .Q(\tms1x00.RAM[95][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4567_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0134_),
    .Q(\tms1x00.RAM[95][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4568_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0135_),
    .Q(\tms1x00.RAM[114][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4569_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0136_),
    .Q(\tms1x00.RAM[114][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4570_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0137_),
    .Q(\tms1x00.RAM[114][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4571_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0138_),
    .Q(\tms1x00.RAM[114][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4572_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0139_),
    .Q(\tms1x00.RAM[113][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4573_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0140_),
    .Q(\tms1x00.RAM[113][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4574_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0141_),
    .Q(\tms1x00.RAM[113][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4575_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0142_),
    .Q(\tms1x00.RAM[113][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4576_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0143_),
    .Q(\tms1x00.RAM[112][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4577_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0144_),
    .Q(\tms1x00.RAM[112][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4578_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0145_),
    .Q(\tms1x00.RAM[112][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4579_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0146_),
    .Q(\tms1x00.RAM[112][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4580_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0147_),
    .Q(\tms1x00.RAM[111][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4581_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0148_),
    .Q(\tms1x00.RAM[111][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4582_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0149_),
    .Q(\tms1x00.RAM[111][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4583_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0150_),
    .Q(\tms1x00.RAM[111][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4584_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0151_),
    .Q(\tms1x00.RAM[110][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4585_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0152_),
    .Q(\tms1x00.RAM[110][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4586_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0153_),
    .Q(\tms1x00.RAM[110][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4587_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0154_),
    .Q(\tms1x00.RAM[110][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4588_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0155_),
    .Q(\tms1x00.RAM[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4589_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0156_),
    .Q(\tms1x00.RAM[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4590_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0157_),
    .Q(\tms1x00.RAM[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4591_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0158_),
    .Q(\tms1x00.RAM[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4592_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0159_),
    .Q(\tms1x00.RAM[108][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4593_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0160_),
    .Q(\tms1x00.RAM[108][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4594_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0161_),
    .Q(\tms1x00.RAM[108][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4595_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0162_),
    .Q(\tms1x00.RAM[108][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4596_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0163_),
    .Q(\tms1x00.RAM[107][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4597_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0164_),
    .Q(\tms1x00.RAM[107][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4598_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0165_),
    .Q(\tms1x00.RAM[107][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4599_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0166_),
    .Q(\tms1x00.RAM[107][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4600_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0167_),
    .Q(\tms1x00.RAM[106][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4601_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0168_),
    .Q(\tms1x00.RAM[106][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4602_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0169_),
    .Q(\tms1x00.RAM[106][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4603_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0170_),
    .Q(\tms1x00.RAM[106][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4604_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0171_),
    .Q(\tms1x00.RAM[105][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4605_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0172_),
    .Q(\tms1x00.RAM[105][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4606_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0173_),
    .Q(\tms1x00.RAM[105][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4607_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0174_),
    .Q(\tms1x00.RAM[105][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4608_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0175_),
    .Q(\tms1x00.RAM[124][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4609_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0176_),
    .Q(\tms1x00.RAM[124][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4610_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0177_),
    .Q(\tms1x00.RAM[124][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4611_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0178_),
    .Q(\tms1x00.RAM[124][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4612_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0179_),
    .Q(\tms1x00.RAM[123][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4613_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0180_),
    .Q(\tms1x00.RAM[123][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4614_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0181_),
    .Q(\tms1x00.RAM[123][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4615_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0182_),
    .Q(\tms1x00.RAM[123][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4616_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0183_),
    .Q(\tms1x00.RAM[122][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4617_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0184_),
    .Q(\tms1x00.RAM[122][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4618_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0185_),
    .Q(\tms1x00.RAM[122][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4619_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0186_),
    .Q(\tms1x00.RAM[122][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4620_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0187_),
    .Q(\tms1x00.RAM[121][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4621_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0188_),
    .Q(\tms1x00.RAM[121][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4622_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0189_),
    .Q(\tms1x00.RAM[121][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4623_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0190_),
    .Q(\tms1x00.RAM[121][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4624_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0191_),
    .Q(\tms1x00.RAM[120][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4625_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0192_),
    .Q(\tms1x00.RAM[120][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4626_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0193_),
    .Q(\tms1x00.RAM[120][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4627_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0194_),
    .Q(\tms1x00.RAM[120][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4628_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0195_),
    .Q(\tms1x00.RAM[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4629_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0196_),
    .Q(\tms1x00.RAM[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4630_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0197_),
    .Q(\tms1x00.RAM[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4631_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0198_),
    .Q(\tms1x00.RAM[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4632_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0199_),
    .Q(\tms1x00.RAM[118][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4633_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0200_),
    .Q(\tms1x00.RAM[118][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4634_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0201_),
    .Q(\tms1x00.RAM[118][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4635_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0202_),
    .Q(\tms1x00.RAM[118][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4636_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0203_),
    .Q(\tms1x00.RAM[117][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4637_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0204_),
    .Q(\tms1x00.RAM[117][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4638_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0205_),
    .Q(\tms1x00.RAM[117][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4639_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0206_),
    .Q(\tms1x00.RAM[117][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4640_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0207_),
    .Q(\tms1x00.RAM[116][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4641_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0208_),
    .Q(\tms1x00.RAM[116][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4642_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0209_),
    .Q(\tms1x00.RAM[116][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4643_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0210_),
    .Q(\tms1x00.RAM[116][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4644_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0211_),
    .Q(\tms1x00.RAM[115][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4645_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0212_),
    .Q(\tms1x00.RAM[115][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4646_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0213_),
    .Q(\tms1x00.RAM[115][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4647_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0214_),
    .Q(\tms1x00.RAM[115][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4648_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0215_),
    .Q(\tms1x00.RAM[126][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4649_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0216_),
    .Q(\tms1x00.RAM[126][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4650_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0217_),
    .Q(\tms1x00.RAM[126][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4651_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0218_),
    .Q(\tms1x00.RAM[126][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4652_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0219_),
    .Q(\tms1x00.RAM[125][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4653_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0220_),
    .Q(\tms1x00.RAM[125][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4654_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0221_),
    .Q(\tms1x00.RAM[125][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4655_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0222_),
    .Q(\tms1x00.RAM[125][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4656_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0223_),
    .Q(\tms1x00.RAM[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4657_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0224_),
    .Q(\tms1x00.RAM[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4658_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0225_),
    .Q(\tms1x00.RAM[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4659_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0226_),
    .Q(\tms1x00.RAM[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4660_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0227_),
    .Q(\tms1x00.RAM[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4661_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0228_),
    .Q(\tms1x00.RAM[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4662_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0229_),
    .Q(\tms1x00.RAM[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4663_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0230_),
    .Q(\tms1x00.RAM[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4664_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0231_),
    .Q(\tms1x00.RAM[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4665_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0232_),
    .Q(\tms1x00.RAM[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4666_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0233_),
    .Q(\tms1x00.RAM[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4667_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0234_),
    .Q(\tms1x00.RAM[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4668_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0235_),
    .Q(\tms1x00.RAM[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4669_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0236_),
    .Q(\tms1x00.RAM[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4670_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0237_),
    .Q(\tms1x00.RAM[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4671_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0238_),
    .Q(\tms1x00.RAM[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4672_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0239_),
    .Q(\tms1x00.RAM[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4673_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0240_),
    .Q(\tms1x00.RAM[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4674_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0241_),
    .Q(\tms1x00.RAM[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4675_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0242_),
    .Q(\tms1x00.RAM[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4676_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0243_),
    .Q(\tms1x00.RAM[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4677_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0244_),
    .Q(\tms1x00.RAM[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4678_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0245_),
    .Q(\tms1x00.RAM[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4679_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0246_),
    .Q(\tms1x00.RAM[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4680_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0247_),
    .Q(\tms1x00.RAM[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4681_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0248_),
    .Q(\tms1x00.RAM[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4682_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0249_),
    .Q(\tms1x00.RAM[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4683_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0250_),
    .Q(\tms1x00.RAM[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4684_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0251_),
    .Q(\tms1x00.RAM[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4685_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0252_),
    .Q(\tms1x00.RAM[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4686_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0253_),
    .Q(\tms1x00.RAM[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4687_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0254_),
    .Q(\tms1x00.RAM[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4688_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0255_),
    .Q(\tms1x00.RAM[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4689_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0256_),
    .Q(\tms1x00.RAM[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4690_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0257_),
    .Q(\tms1x00.RAM[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4691_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0258_),
    .Q(\tms1x00.RAM[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4692_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0259_),
    .Q(\tms1x00.RAM[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4693_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0260_),
    .Q(\tms1x00.RAM[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4694_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0261_),
    .Q(\tms1x00.RAM[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4695_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0262_),
    .Q(\tms1x00.RAM[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4696_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0263_),
    .Q(\tms1x00.RAM[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4697_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0264_),
    .Q(\tms1x00.RAM[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4698_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0265_),
    .Q(\tms1x00.RAM[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4699_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0266_),
    .Q(\tms1x00.RAM[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4700_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0267_),
    .Q(\tms1x00.RAM[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4701_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0268_),
    .Q(\tms1x00.RAM[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4702_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0269_),
    .Q(\tms1x00.RAM[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4703_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0270_),
    .Q(\tms1x00.RAM[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4704_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0271_),
    .Q(\tms1x00.RAM[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4705_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0272_),
    .Q(\tms1x00.RAM[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4706_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0273_),
    .Q(\tms1x00.RAM[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4707_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0274_),
    .Q(\tms1x00.RAM[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4708_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0275_),
    .Q(\tms1x00.RAM[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4709_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0276_),
    .Q(\tms1x00.RAM[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4710_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0277_),
    .Q(\tms1x00.RAM[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4711_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0278_),
    .Q(\tms1x00.RAM[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4712_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0279_),
    .Q(\tms1x00.RAM[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4713_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0280_),
    .Q(\tms1x00.RAM[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4714_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0281_),
    .Q(\tms1x00.RAM[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4715_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0282_),
    .Q(\tms1x00.RAM[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4716_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0283_),
    .Q(\tms1x00.RAM[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4717_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0284_),
    .Q(\tms1x00.RAM[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4718_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0285_),
    .Q(\tms1x00.RAM[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4719_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0286_),
    .Q(\tms1x00.RAM[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _4720_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0042_),
    .Q(_0035_));
 sky130_fd_sc_hd__dfxtp_1 _4721_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0043_),
    .Q(_0036_));
 sky130_fd_sc_hd__dfxtp_1 _4722_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0044_),
    .Q(_0037_));
 sky130_fd_sc_hd__dfxtp_4 _4723_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0045_),
    .Q(_0038_));
 sky130_fd_sc_hd__dfxtp_4 _4724_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0046_),
    .Q(_0039_));
 sky130_fd_sc_hd__dfxtp_4 _4725_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0047_),
    .Q(_0040_));
 sky130_fd_sc_hd__dfxtp_2 _4726_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0048_),
    .Q(_0041_));
 sky130_fd_sc_hd__dfxtp_1 _4727_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0287_),
    .Q(\tms1x00.RAM[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4728_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0288_),
    .Q(\tms1x00.RAM[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4729_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0289_),
    .Q(\tms1x00.RAM[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4730_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0290_),
    .Q(\tms1x00.RAM[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4731_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0291_),
    .Q(\tms1x00.RAM[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4732_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0292_),
    .Q(\tms1x00.RAM[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4733_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0293_),
    .Q(\tms1x00.RAM[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4734_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0294_),
    .Q(\tms1x00.RAM[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4735_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0295_),
    .Q(\tms1x00.RAM[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4736_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0296_),
    .Q(\tms1x00.RAM[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4737_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0297_),
    .Q(\tms1x00.RAM[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4738_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0298_),
    .Q(\tms1x00.RAM[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4739_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0299_),
    .Q(\tms1x00.RAM[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4740_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0300_),
    .Q(\tms1x00.RAM[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4741_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0301_),
    .Q(\tms1x00.RAM[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4742_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0302_),
    .Q(\tms1x00.RAM[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4743_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0303_),
    .Q(\tms1x00.RAM[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4744_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0304_),
    .Q(\tms1x00.RAM[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4745_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0305_),
    .Q(\tms1x00.RAM[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4746_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0306_),
    .Q(\tms1x00.RAM[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4747_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0307_),
    .Q(\tms1x00.RAM[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4748_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0308_),
    .Q(\tms1x00.RAM[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4749_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0309_),
    .Q(\tms1x00.RAM[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4750_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0310_),
    .Q(\tms1x00.RAM[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4751_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0311_),
    .Q(\tms1x00.RAM[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4752_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0312_),
    .Q(\tms1x00.RAM[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4753_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0313_),
    .Q(\tms1x00.RAM[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4754_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0314_),
    .Q(\tms1x00.RAM[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4755_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0315_),
    .Q(\tms1x00.RAM[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4756_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0316_),
    .Q(\tms1x00.RAM[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4757_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0317_),
    .Q(\tms1x00.RAM[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4758_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0318_),
    .Q(\tms1x00.RAM[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4759_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0319_),
    .Q(\tms1x00.RAM[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4760_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0320_),
    .Q(\tms1x00.RAM[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4761_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0321_),
    .Q(\tms1x00.RAM[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4762_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0322_),
    .Q(\tms1x00.RAM[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4763_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0323_),
    .Q(\tms1x00.RAM[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4764_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0324_),
    .Q(\tms1x00.RAM[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4765_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0325_),
    .Q(\tms1x00.RAM[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4766_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0326_),
    .Q(\tms1x00.RAM[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4767_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0327_),
    .Q(\tms1x00.RAM[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4768_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0328_),
    .Q(\tms1x00.RAM[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4769_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0329_),
    .Q(\tms1x00.RAM[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4770_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0330_),
    .Q(\tms1x00.RAM[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4771_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0331_),
    .Q(\tms1x00.RAM[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4772_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0332_),
    .Q(\tms1x00.RAM[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4773_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0333_),
    .Q(\tms1x00.RAM[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4774_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0334_),
    .Q(\tms1x00.RAM[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4775_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0335_),
    .Q(\tms1x00.RAM[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4776_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0336_),
    .Q(\tms1x00.RAM[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4777_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0337_),
    .Q(\tms1x00.RAM[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4778_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0338_),
    .Q(\tms1x00.RAM[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4779_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0339_),
    .Q(\tms1x00.RAM[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4780_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0340_),
    .Q(\tms1x00.RAM[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4781_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0341_),
    .Q(\tms1x00.RAM[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4782_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0342_),
    .Q(\tms1x00.RAM[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4783_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0343_),
    .Q(\tms1x00.RAM[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4784_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0344_),
    .Q(\tms1x00.RAM[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4785_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0345_),
    .Q(\tms1x00.RAM[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4786_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0346_),
    .Q(\tms1x00.RAM[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4787_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0347_),
    .Q(\tms1x00.RAM[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4788_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0348_),
    .Q(\tms1x00.RAM[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4789_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0349_),
    .Q(\tms1x00.RAM[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4790_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0350_),
    .Q(\tms1x00.RAM[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4791_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0351_),
    .Q(\tms1x00.RAM[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4792_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0352_),
    .Q(\tms1x00.RAM[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4793_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0353_),
    .Q(\tms1x00.RAM[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4794_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0354_),
    .Q(\tms1x00.RAM[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4795_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0355_),
    .Q(\tms1x00.RAM[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4796_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0356_),
    .Q(\tms1x00.RAM[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4797_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0357_),
    .Q(\tms1x00.RAM[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4798_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0358_),
    .Q(\tms1x00.RAM[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4799_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0359_),
    .Q(\tms1x00.RAM[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4800_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0360_),
    .Q(\tms1x00.RAM[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4801_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0361_),
    .Q(\tms1x00.RAM[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4802_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0362_),
    .Q(\tms1x00.RAM[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4803_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0363_),
    .Q(\tms1x00.RAM[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4804_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0364_),
    .Q(\tms1x00.RAM[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4805_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0365_),
    .Q(\tms1x00.RAM[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4806_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0366_),
    .Q(\tms1x00.RAM[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4807_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0367_),
    .Q(\tms1x00.RAM[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4808_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0368_),
    .Q(\tms1x00.RAM[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4809_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0369_),
    .Q(\tms1x00.RAM[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4810_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0370_),
    .Q(\tms1x00.RAM[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4811_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0371_),
    .Q(\tms1x00.RAM[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4812_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0372_),
    .Q(\tms1x00.RAM[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4813_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0373_),
    .Q(\tms1x00.RAM[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4814_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0374_),
    .Q(\tms1x00.RAM[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4815_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0375_),
    .Q(\tms1x00.RAM[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4816_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0376_),
    .Q(\tms1x00.RAM[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4817_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0377_),
    .Q(\tms1x00.RAM[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4818_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0378_),
    .Q(\tms1x00.RAM[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4819_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0379_),
    .Q(\tms1x00.RAM[67][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4820_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0380_),
    .Q(\tms1x00.RAM[67][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4821_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0381_),
    .Q(\tms1x00.RAM[67][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4822_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0382_),
    .Q(\tms1x00.RAM[67][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4823_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0383_),
    .Q(\tms1x00.RAM[66][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4824_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0384_),
    .Q(\tms1x00.RAM[66][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4825_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0385_),
    .Q(\tms1x00.RAM[66][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4826_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0386_),
    .Q(\tms1x00.RAM[66][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4827_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0387_),
    .Q(\tms1x00.RAM[65][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4828_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0388_),
    .Q(\tms1x00.RAM[65][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4829_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0389_),
    .Q(\tms1x00.RAM[65][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4830_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0390_),
    .Q(\tms1x00.RAM[65][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4831_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0391_),
    .Q(\tms1x00.RAM[64][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4832_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0392_),
    .Q(\tms1x00.RAM[64][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4833_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0393_),
    .Q(\tms1x00.RAM[64][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4834_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0394_),
    .Q(\tms1x00.RAM[64][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4835_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0395_),
    .Q(\tms1x00.RAM[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4836_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0396_),
    .Q(\tms1x00.RAM[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4837_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0397_),
    .Q(\tms1x00.RAM[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4838_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0398_),
    .Q(\tms1x00.RAM[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4839_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0399_),
    .Q(\tms1x00.RAM[71][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4840_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0400_),
    .Q(\tms1x00.RAM[71][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4841_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0401_),
    .Q(\tms1x00.RAM[71][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4842_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0402_),
    .Q(\tms1x00.RAM[71][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4843_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0403_),
    .Q(\tms1x00.RAM[70][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4844_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0404_),
    .Q(\tms1x00.RAM[70][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4845_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0405_),
    .Q(\tms1x00.RAM[70][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4846_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0406_),
    .Q(\tms1x00.RAM[70][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4847_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0407_),
    .Q(\tms1x00.RAM[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4848_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0408_),
    .Q(\tms1x00.RAM[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4849_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0409_),
    .Q(\tms1x00.RAM[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4850_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0410_),
    .Q(\tms1x00.RAM[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4851_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0411_),
    .Q(\tms1x00.RAM[68][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4852_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0412_),
    .Q(\tms1x00.RAM[68][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4853_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0413_),
    .Q(\tms1x00.RAM[68][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4854_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0414_),
    .Q(\tms1x00.RAM[68][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4855_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0415_),
    .Q(\tms1x00.RAM[76][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4856_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0416_),
    .Q(\tms1x00.RAM[76][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4857_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0417_),
    .Q(\tms1x00.RAM[76][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4858_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0418_),
    .Q(\tms1x00.RAM[76][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4859_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0419_),
    .Q(\tms1x00.RAM[75][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4860_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0420_),
    .Q(\tms1x00.RAM[75][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4861_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0421_),
    .Q(\tms1x00.RAM[75][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4862_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0422_),
    .Q(\tms1x00.RAM[75][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4863_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0423_),
    .Q(\tms1x00.RAM[74][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4864_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0424_),
    .Q(\tms1x00.RAM[74][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4865_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0425_),
    .Q(\tms1x00.RAM[74][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4866_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0426_),
    .Q(\tms1x00.RAM[74][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4867_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0427_),
    .Q(\tms1x00.RAM[73][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4868_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0428_),
    .Q(\tms1x00.RAM[73][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4869_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0429_),
    .Q(\tms1x00.RAM[73][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4870_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0430_),
    .Q(\tms1x00.RAM[73][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4871_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0431_),
    .Q(\tms1x00.RAM[72][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4872_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0432_),
    .Q(\tms1x00.RAM[72][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4873_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0433_),
    .Q(\tms1x00.RAM[72][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4874_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0434_),
    .Q(\tms1x00.RAM[72][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4875_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0435_),
    .Q(\tms1x00.RAM[80][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4876_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0436_),
    .Q(\tms1x00.RAM[80][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4877_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0437_),
    .Q(\tms1x00.RAM[80][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4878_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0438_),
    .Q(\tms1x00.RAM[80][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4879_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0439_),
    .Q(\tms1x00.RAM[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4880_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0440_),
    .Q(\tms1x00.RAM[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4881_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0441_),
    .Q(\tms1x00.RAM[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4882_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0442_),
    .Q(\tms1x00.RAM[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4883_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0443_),
    .Q(\tms1x00.RAM[78][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4884_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0444_),
    .Q(\tms1x00.RAM[78][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4885_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0445_),
    .Q(\tms1x00.RAM[78][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4886_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0446_),
    .Q(\tms1x00.RAM[78][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4887_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0447_),
    .Q(\tms1x00.RAM[77][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4888_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0448_),
    .Q(\tms1x00.RAM[77][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4889_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0449_),
    .Q(\tms1x00.RAM[77][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4890_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0450_),
    .Q(\tms1x00.RAM[77][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4891_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0451_),
    .Q(\tms1x00.RAM[85][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4892_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0452_),
    .Q(\tms1x00.RAM[85][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4893_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0453_),
    .Q(\tms1x00.RAM[85][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4894_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0454_),
    .Q(\tms1x00.RAM[85][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4895_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0455_),
    .Q(\tms1x00.RAM[84][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4896_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0456_),
    .Q(\tms1x00.RAM[84][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4897_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0457_),
    .Q(\tms1x00.RAM[84][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4898_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0458_),
    .Q(\tms1x00.RAM[84][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4899_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0459_),
    .Q(\tms1x00.RAM[83][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4900_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0460_),
    .Q(\tms1x00.RAM[83][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4901_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0461_),
    .Q(\tms1x00.RAM[83][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4902_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0462_),
    .Q(\tms1x00.RAM[83][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4903_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0463_),
    .Q(\tms1x00.RAM[82][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4904_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0464_),
    .Q(\tms1x00.RAM[82][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4905_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0465_),
    .Q(\tms1x00.RAM[82][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4906_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0466_),
    .Q(\tms1x00.RAM[82][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4907_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0467_),
    .Q(\tms1x00.RAM[81][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4908_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0468_),
    .Q(\tms1x00.RAM[81][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4909_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0469_),
    .Q(\tms1x00.RAM[81][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4910_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0470_),
    .Q(\tms1x00.RAM[81][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4911_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0471_),
    .Q(\tms1x00.RAM[86][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4912_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0472_),
    .Q(\tms1x00.RAM[86][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4913_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0473_),
    .Q(\tms1x00.RAM[86][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4914_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0474_),
    .Q(\tms1x00.RAM[86][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4915_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0475_),
    .Q(\tms1x00.RAM[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4916_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0476_),
    .Q(\tms1x00.RAM[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4917_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0477_),
    .Q(\tms1x00.RAM[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4918_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0478_),
    .Q(\tms1x00.RAM[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4919_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0479_),
    .Q(\tms1x00.RAM[88][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4920_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0480_),
    .Q(\tms1x00.RAM[88][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4921_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0481_),
    .Q(\tms1x00.RAM[88][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4922_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0482_),
    .Q(\tms1x00.RAM[88][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4923_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0483_),
    .Q(\tms1x00.RAM[87][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4924_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0484_),
    .Q(\tms1x00.RAM[87][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4925_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0485_),
    .Q(\tms1x00.RAM[87][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4926_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0486_),
    .Q(\tms1x00.RAM[87][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4927_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0487_),
    .Q(\tms1x00.RAM[94][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4928_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0488_),
    .Q(\tms1x00.RAM[94][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4929_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0489_),
    .Q(\tms1x00.RAM[94][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4930_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0490_),
    .Q(\tms1x00.RAM[94][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4931_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0491_),
    .Q(\tms1x00.RAM[93][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4932_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0492_),
    .Q(\tms1x00.RAM[93][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4933_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0493_),
    .Q(\tms1x00.RAM[93][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4934_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0494_),
    .Q(\tms1x00.RAM[93][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4935_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0495_),
    .Q(\tms1x00.RAM[92][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4936_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0496_),
    .Q(\tms1x00.RAM[92][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4937_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0497_),
    .Q(\tms1x00.RAM[92][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4938_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0498_),
    .Q(\tms1x00.RAM[92][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4939_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0499_),
    .Q(\tms1x00.RAM[91][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4940_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0500_),
    .Q(\tms1x00.RAM[91][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4941_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0501_),
    .Q(\tms1x00.RAM[91][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4942_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0502_),
    .Q(\tms1x00.RAM[91][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4943_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0503_),
    .Q(\tms1x00.RAM[90][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4944_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0504_),
    .Q(\tms1x00.RAM[90][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4945_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0505_),
    .Q(\tms1x00.RAM[90][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4946_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0506_),
    .Q(\tms1x00.RAM[90][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4947_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0507_),
    .Q(\tms1x00.RAM[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4948_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0508_),
    .Q(\tms1x00.RAM[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4949_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0509_),
    .Q(\tms1x00.RAM[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4950_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0510_),
    .Q(\tms1x00.RAM[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4951_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0511_),
    .Q(\tms1x00.ram_addr_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4952_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0512_),
    .Q(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4953_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0513_),
    .Q(\tms1x00.ram_addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4954_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0514_),
    .Q(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_4 _4955_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0515_),
    .Q(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_4 _4956_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0516_),
    .Q(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_4 _4957_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0517_),
    .Q(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4958_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0518_),
    .Q(\tms1x00.wb_step_state ));
 sky130_fd_sc_hd__dfxtp_4 _4959_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0519_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_2 _4960_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0520_),
    .Q(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4961_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0521_),
    .Q(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4962_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0522_),
    .Q(\tms1x00.ins_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4963_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0523_),
    .Q(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4964_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0524_),
    .Q(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4965_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0525_),
    .Q(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__dfxtp_2 _4966_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0526_),
    .Q(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4967_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0527_),
    .Q(\tms1x00.ins_in[7] ));
 sky130_fd_sc_hd__dfxtp_2 _4968_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0528_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_4 _4969_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0529_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_4 _4970_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0530_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _4971_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(\tms1x00.K_in[0] ),
    .Q(\tms1x00.K_latch[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4972_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(\tms1x00.K_in[1] ),
    .Q(\tms1x00.K_latch[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4973_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\tms1x00.K_in[2] ),
    .Q(\tms1x00.K_latch[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4974_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(\tms1x00.K_in[3] ),
    .Q(\tms1x00.K_latch[3] ));
 sky130_fd_sc_hd__dfxtp_4 _4975_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0531_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_4 _4976_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0532_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_4 _4977_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0533_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_4 _4978_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0534_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_2 _4979_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0535_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_4 _4980_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0536_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_4 _4981_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0537_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_4 _4982_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0538_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_4 _4983_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0539_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_4 _4984_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0540_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_4 _4985_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0541_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_4 _4986_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0542_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_4 _4987_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0543_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_4 _4988_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0544_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_4 _4989_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0545_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_2 _4990_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0546_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_2 _4991_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0547_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_2 _4992_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0548_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_2 _4993_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0549_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_2 _4994_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0550_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_2 _4995_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0551_),
    .Q(\tms1x00.CL ));
 sky130_fd_sc_hd__dfxtp_1 _4996_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0552_),
    .Q(\tms1x00.status ));
 sky130_fd_sc_hd__dfxtp_1 _4997_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0553_),
    .Q(\tms1x00.SR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4998_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0554_),
    .Q(\tms1x00.SR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4999_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0555_),
    .Q(\tms1x00.SR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5000_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0556_),
    .Q(\tms1x00.SR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5001_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0557_),
    .Q(\tms1x00.SR[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5002_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0558_),
    .Q(\tms1x00.SR[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5003_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0559_),
    .Q(\tms1x00.PB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5004_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0560_),
    .Q(\tms1x00.PB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5005_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0561_),
    .Q(\tms1x00.PB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5006_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0562_),
    .Q(\tms1x00.PB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5007_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0563_),
    .Q(\tms1x00.PA[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5008_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0564_),
    .Q(\tms1x00.PA[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5009_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0565_),
    .Q(\tms1x00.PA[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5010_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0566_),
    .Q(\tms1x00.PA[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5011_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0567_),
    .Q(\tms1x00.P[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5012_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0568_),
    .Q(\tms1x00.P[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5013_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0569_),
    .Q(\tms1x00.P[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5014_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0570_),
    .Q(\tms1x00.P[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5015_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0571_),
    .Q(\tms1x00.PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5016_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0572_),
    .Q(\tms1x00.PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5017_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0573_),
    .Q(\tms1x00.PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5018_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0574_),
    .Q(\tms1x00.PC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5019_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0575_),
    .Q(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5020_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0576_),
    .Q(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__dfxtp_2 _5021_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0577_),
    .Q(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__dfxtp_2 _5022_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0578_),
    .Q(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5023_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0579_),
    .Q(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5024_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0580_),
    .Q(\tms1x00.Y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5025_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0581_),
    .Q(\tms1x00.X[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5026_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0582_),
    .Q(\tms1x00.X[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5027_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0583_),
    .Q(\tms1x00.X[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5028_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0584_),
    .Q(\tms1x00.N[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5029_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0585_),
    .Q(\tms1x00.N[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5030_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0586_),
    .Q(\tms1x00.N[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5031_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0587_),
    .Q(\tms1x00.N[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5032_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0588_),
    .Q(\tms1x00.A[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5033_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0589_),
    .Q(\tms1x00.A[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5034_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0590_),
    .Q(\tms1x00.A[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5035_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0591_),
    .Q(\tms1x00.A[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5036_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0592_),
    .Q(\tms1x00.RAM[119][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5037_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0593_),
    .Q(\tms1x00.RAM[119][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5038_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0594_),
    .Q(\tms1x00.RAM[119][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5039_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0595_),
    .Q(\tms1x00.RAM[119][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5040_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0596_),
    .Q(\tms1x00.RAM[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5041_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0597_),
    .Q(\tms1x00.RAM[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5042_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0598_),
    .Q(\tms1x00.RAM[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5043_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0599_),
    .Q(\tms1x00.RAM[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5044_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0600_),
    .Q(\tms1x00.RAM[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5045_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0601_),
    .Q(\tms1x00.RAM[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5046_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0602_),
    .Q(\tms1x00.RAM[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5047_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0603_),
    .Q(\tms1x00.RAM[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5048_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0604_),
    .Q(\tms1x00.RAM[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5049_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0605_),
    .Q(\tms1x00.RAM[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5050_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0606_),
    .Q(\tms1x00.RAM[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5051_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0607_),
    .Q(\tms1x00.RAM[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5052_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0608_),
    .Q(\tms1x00.RAM[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5053_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0609_),
    .Q(\tms1x00.RAM[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5054_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0610_),
    .Q(\tms1x00.RAM[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5055_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0611_),
    .Q(\tms1x00.RAM[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5056_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0612_),
    .Q(\tms1x00.RAM[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5057_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0613_),
    .Q(\tms1x00.RAM[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5058_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0614_),
    .Q(\tms1x00.RAM[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5059_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0615_),
    .Q(\tms1x00.RAM[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5060_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0616_),
    .Q(\tms1x00.RAM[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5061_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0617_),
    .Q(\tms1x00.RAM[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5062_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0618_),
    .Q(\tms1x00.RAM[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5063_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0619_),
    .Q(\tms1x00.RAM[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5064_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0620_),
    .Q(\tms1x00.RAM[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5065_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0621_),
    .Q(\tms1x00.RAM[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5066_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0622_),
    .Q(\tms1x00.RAM[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5067_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0623_),
    .Q(\tms1x00.RAM[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5068_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0624_),
    .Q(\tms1x00.RAM[127][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5069_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0625_),
    .Q(\tms1x00.RAM[127][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5070_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0626_),
    .Q(\tms1x00.RAM[127][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5071_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0627_),
    .Q(\tms1x00.RAM[127][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5072_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0628_),
    .Q(\tms1x00.RAM[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5073_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0629_),
    .Q(\tms1x00.RAM[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5074_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0630_),
    .Q(\tms1x00.RAM[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5075_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0631_),
    .Q(\tms1x00.RAM[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5076_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0632_),
    .Q(\tms1x00.RAM[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5077_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0633_),
    .Q(\tms1x00.RAM[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5078_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0634_),
    .Q(\tms1x00.RAM[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5079_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0635_),
    .Q(\tms1x00.RAM[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5080_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0636_),
    .Q(\tms1x00.RAM[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5081_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0637_),
    .Q(\tms1x00.RAM[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5082_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0638_),
    .Q(\tms1x00.RAM[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5083_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0639_),
    .Q(\tms1x00.RAM[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5084_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0640_),
    .Q(\tms1x00.RAM[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5085_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0641_),
    .Q(\tms1x00.RAM[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5086_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0642_),
    .Q(\tms1x00.RAM[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5087_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0643_),
    .Q(\tms1x00.RAM[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5088_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0644_),
    .Q(\tms1x00.RAM[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5089_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0645_),
    .Q(\tms1x00.RAM[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5090_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0646_),
    .Q(\tms1x00.RAM[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5091_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0647_),
    .Q(\tms1x00.RAM[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _5092_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0648_),
    .Q(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _5093_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0649_),
    .Q(\tms1x00.rom_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5094_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0650_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _5095_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0651_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _5096_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0652_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _5097_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0653_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _5098_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0654_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_1 _5099_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0655_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_1 _5100_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0656_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_1 _5101_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0657_),
    .Q(net105));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_195 (.HI(net195));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_196 (.HI(net196));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_197 (.HI(net197));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_198 (.HI(net198));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_199 (.HI(net199));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_200 (.HI(net200));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_201 (.HI(net201));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_202 (.HI(net202));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_203 (.HI(net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_166 (.LO(net166));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_167 (.LO(net167));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_168 (.LO(net168));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_169 (.LO(net169));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_170 (.LO(net170));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_171 (.LO(net171));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_172 (.LO(net172));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_173 (.LO(net173));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_174 (.LO(net174));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_175 (.LO(net175));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_176 (.LO(net176));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_177 (.LO(net177));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_178 (.LO(net178));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_179 (.LO(net179));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_180 (.LO(net180));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_181 (.LO(net181));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_182 (.LO(net182));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_183 (.LO(net183));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_184 (.LO(net184));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_190 (.LO(net190));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_191 (.LO(net191));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_192 (.LO(net192));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_193 (.LO(net193));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_194 (.HI(net194));
 sky130_fd_sc_hd__clkbuf_1 _5153_ (.A(net53),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 _5154_ (.A(net54),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 _5155_ (.A(net55),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 _5156_ (.A(net56),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 _5157_ (.A(net57),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 _5158_ (.A(net58),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 _5159_ (.A(net59),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 _5160_ (.A(net60),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 _5161_ (.A(net50),
    .X(net115));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[5]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[6]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[7]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[8]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[9]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(oram_value[0]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(oram_value[10]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(oram_value[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(oram_value[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(oram_value[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(oram_value[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(oram_value[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(oram_value[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(oram_value[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(oram_value[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(oram_value[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(ram_val[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(ram_val[10]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(ram_val[11]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(ram_val[12]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(ram_val[13]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(ram_val[14]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(ram_val[15]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(ram_val[16]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(ram_val[17]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(ram_val[18]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(ram_val[19]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(ram_val[1]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(ram_val[20]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(ram_val[21]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(ram_val[22]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(ram_val[23]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(ram_val[24]),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(ram_val[25]),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(ram_val[26]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(ram_val[27]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(ram_val[28]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(ram_val[29]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(ram_val[2]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(ram_val[30]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(ram_val[31]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(ram_val[3]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(ram_val[4]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(ram_val[5]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(ram_val[6]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(ram_val[7]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(ram_val[8]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(ram_val[9]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(wb_rst_i),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(wbs_adr_i[10]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(wbs_adr_i[16]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(wbs_adr_i[23]),
    .X(net52));
 sky130_fd_sc_hd__dlymetal6s2s_1 input53 (.A(wbs_adr_i[2]),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 input54 (.A(wbs_adr_i[3]),
    .X(net54));
 sky130_fd_sc_hd__dlymetal6s2s_1 input55 (.A(wbs_adr_i[4]),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(wbs_adr_i[5]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(wbs_adr_i[6]),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(wbs_adr_i[7]),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 input59 (.A(wbs_adr_i[8]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(wbs_adr_i[9]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(wbs_cyc_i),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(wbs_dat_i[0]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(wbs_dat_i[10]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(wbs_dat_i[11]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(wbs_dat_i[1]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(wbs_dat_i[2]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(wbs_dat_i[3]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(wbs_dat_i[8]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(wbs_dat_i[9]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(wbs_stb_i),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(wbs_we_i),
    .X(net71));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(io_out[36]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(io_out[37]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(oram_addr[0]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(oram_addr[1]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(oram_addr[2]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(oram_addr[3]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(oram_addr[4]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(oram_addr[5]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(oram_addr[6]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(oram_addr[7]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(oram_csb));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(ram_adrb[0]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(ram_adrb[1]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(ram_adrb[2]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(ram_adrb[3]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(ram_adrb[4]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(ram_adrb[5]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(ram_adrb[6]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(ram_adrb[7]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(ram_adrb[8]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(ram_csb));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(ram_web));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(net77),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net97),
    .X(net152));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_153 (.LO(net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_wb_clk_i (.A(clknet_1_0_0_wb_clk_i),
    .X(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_wb_clk_i (.A(clknet_1_0_0_wb_clk_i),
    .X(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_wb_clk_i (.A(clknet_1_1_0_wb_clk_i),
    .X(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_wb_clk_i (.A(clknet_1_1_0_wb_clk_i),
    .X(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(feedback_delay),
    .X(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__A0 (.DIODE(\K_override[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__A1 (.DIODE(\K_override[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__A0 (.DIODE(\K_override[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__A1 (.DIODE(\K_override[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__A0 (.DIODE(\K_override[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__A1 (.DIODE(\K_override[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__A0 (.DIODE(\K_override[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__A1 (.DIODE(\K_override[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__A (.DIODE(_0037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__A (.DIODE(_0037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__B1 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__B1 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__B1 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__A (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__A (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__A (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2857__C1 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__C1 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2714__C1 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__A1 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__B1 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__C1 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__A (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__A (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2858__C1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__B1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__A1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__A1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__C1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__C1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__A1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__C1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__A (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2860__A1 (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__B1 (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__C1 (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__B1 (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__A (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A2 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2314__A2 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2313__A2 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__A2 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__A (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__B (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2286__A (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2300__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2288__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__B (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__B (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__B (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__B (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__B (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__B (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2314__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2313__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__C (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__A1 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__A1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__B2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A0 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__A0 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__B2 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A1 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A1 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__A1 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A1 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A1 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A1 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__A1 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__A (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A1 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A1 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__A1 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A1 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__A0 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2393__A1 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__A0 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__B_N (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__A1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__A1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__B (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__A2 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__B (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__A1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__D (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__B (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__B (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__B (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__B (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A3 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__A3 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2390__A (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__C1 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__C1 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__C1 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__C1 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__B1 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__B1 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__B (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2393__C1 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2656__B1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__B1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__B1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__A (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2856__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2758__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2713__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2704__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__C1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__A (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2825__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__C1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__C1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__S0 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__S0 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__S0 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__S0 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__S0 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__S0 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__S0 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__S0 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__A (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__A (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2835__S (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2811__S0 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2805__S0 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2643__S0 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__S0 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__S0 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__S0 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__S0 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__S0 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__S0 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__S1 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__S1 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__S1 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__S1 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__S1 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__S1 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__S1 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__A (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__A (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2805__S1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2754__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2643__S1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__S1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__S1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__S1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__S1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__S1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__S1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__S1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__S0 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__S0 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__S0 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__S0 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__S0 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__S (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__S (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__A (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__S0 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__S0 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__S0 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__S0 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__S (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__S0 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__S0 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2641__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2426__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2854__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2797__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2745__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__A1 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2711__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__S (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__S (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__S1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__S1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__S1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__S1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__S1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2417__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2412__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__S1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__S1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__S1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__A (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__B1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__B1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__A (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__B1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__B1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__A (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2816__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__A (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__B1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2416__A (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__A (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2836__B2 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__A1 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__A1 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__B2 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__A1 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__B2 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__A1 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__B2 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__A1 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__A1 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__S0 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__A (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2607__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2439__A (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2420__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__C1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__A (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__C1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__A (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__C1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__A (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__A (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__B1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2845__B1 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2811__S1 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__B1 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2628__B1 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__S1 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__S1 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__S1 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__S1 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__S1 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__S1 (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__A1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__A1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__B2 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__B2 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__A1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2502__A (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__A1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__B2 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__B2 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__C1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__C1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2824__B1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2793__C1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__C1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__C1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__B1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2499__B1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__C1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__C1 (.DIODE(_0795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__C1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2705__C1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2657__C1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__C1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__C1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__C1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2430__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2858__A1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2825__C1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2813__C1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__C1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__C1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__C1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__C1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__C1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__C1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__C1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__A2 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2852__B1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__B1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__B1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__B1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__B1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__B1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2642__C1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__B1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__B1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__A (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__C1 (.DIODE(_0801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__C1 (.DIODE(_0801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__A1 (.DIODE(_0801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__B1 (.DIODE(_0801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2694__A1 (.DIODE(_0801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2679__C1 (.DIODE(_0801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__A1 (.DIODE(_0801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__A1 (.DIODE(_0801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__A1 (.DIODE(_0801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__A1 (.DIODE(_0801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2852__A1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2804__A (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2758__A1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__A1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2704__A1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__B2 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__A (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__A (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__S (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__A (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__S0 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2803__S0 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__S0 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__S0 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__S0 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__S0 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__B_N (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2475__B_N (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__S0 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__S1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2803__S1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2790__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__S1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__S1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__S1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__S1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__S1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__A (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__S1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2832__S0 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__S0 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__S0 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__S0 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2626__B_N (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__A1 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__B_N (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__S (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__A1 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__B_N (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2808__B1 (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__A (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2618__A (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__S1 (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__A (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__B1 (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__S1 (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__S1 (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__A (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__B1 (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__S0 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__S0 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__S0 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__S0 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__S0 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__S0 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__S0 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__S0 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__S0 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__A (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2735__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__S0 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2847__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2792__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__A1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__A1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2702__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2654__C1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__A1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2645__A (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__B1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__A (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__B1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__B1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__A (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__B1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__A (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2856__A1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__C1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__B1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2713__A1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__A1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2691__B1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__B1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2642__A1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__C1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__C1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2838__A (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__A1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2794__A (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__B1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2694__B1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__A1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__B1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__B1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__B1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__B1 (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__C1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2831__C1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__C1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__C1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__C1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__C1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__C1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__C1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__C1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__C1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__A1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2821__B1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__A1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__A1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__C1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2722__B1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__C1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__A1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__C1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__A1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__S (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2791__S (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__S (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__S (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__S (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__S0 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__S0 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__S0 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__S0 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__S0 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__S1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__S1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__S1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__S1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__S1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__S1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__S1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__S1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__S1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__S1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2851__S0 (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__S (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2800__S0 (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__S0 (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__S0 (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__A1 (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__B_N (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__S0 (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__A (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A1 (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__A (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2656__A1 (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__A1 (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__S (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__A1 (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__A (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__A (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__A1 (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__A (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__A1 (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__B1 (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__A (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__B1 (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2822__A1 (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__A1 (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__B2 (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2723__A1 (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2691__A1 (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__B2 (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__A1 (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__A1 (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__B2 (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__A1 (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2823__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__A1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__B_N (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__S (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2823__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__A (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__A1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2836__C1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2792__C1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2741__A (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__A1 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2831__B2 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2818__S (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__B2 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__S (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__A (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__S (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__S (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__B2 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2499__A1 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2834__A1 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2833__B_N (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__S0 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2809__S (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2790__A1 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__B_N (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__S (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2754__A1 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__S (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__S (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__A2 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__A2 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__B (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__A2 (.DIODE(_0894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__B (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__B2 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__A (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2551__A (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3097__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2879__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__A0 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A0 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A0 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__A0 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2998__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2871__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3061__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2870__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__C (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__C (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__A (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__A (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__A (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__B (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__S0 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__S0 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__S0 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__S0 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2742__S0 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2710__S0 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2695__S0 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__S0 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__S0 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__S0 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__S1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2849__S1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2796__S1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__S1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__S1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2742__S1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__S1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2695__S1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__S1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__S1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2843__S1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2839__S1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2832__S1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2827__A (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__S1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2788__S1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__S1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__S1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__S1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__A1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2849__S0 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2796__S0 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__S0 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__S0 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__S0 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__S0 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2681__A (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__A1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__B_N (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__S (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2613__A2 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2851__S1 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2834__B1 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2800__S1 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__S1 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__S1 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2710__S1 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__S1 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__S1 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__S1 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__S1 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__B1 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__B1 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A (.DIODE(_0980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__A1 (.DIODE(_0980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__B1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2845__A1 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__B_N (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2820__S (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__S0 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2816__S0 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2753__B_N (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2721__S (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__A1 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__B_N (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2628__A1 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__B1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2850__A (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2847__C1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2801__A (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__C1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__A1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__B1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__A (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2702__C1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__C1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__A2 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__A2 (.DIODE(_1016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2656__A2 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__A2 (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3035__A (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__A (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__A (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__A (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2887__A (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__A (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A0 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A0 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__A0 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__A0 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3012__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2873__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2821__A1 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__S1 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__A (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__A (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__B1 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2722__A1 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__A (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2685__B1 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2677__S1 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2673__A (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2819__S (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__S0 (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__S (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__A1 (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__B_N (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2720__S (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2686__S (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2685__A1 (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__B_N (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2677__S0 (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__A1 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2824__A1 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__A1 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2793__A1 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__B2 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__B2 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__A1 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__B2 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__A (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2679__B2 (.DIODE(_1044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2716__A2 (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2843__S0 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2839__S0 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2808__A1 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2807__B_N (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__S0 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2788__S0 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__S0 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__S0 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__S0 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__S0 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2702__B1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__A2 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__A (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__A1 (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__A2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__B1 (.DIODE(_1097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A2 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__B (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__A2 (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__A (.DIODE(_1131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__A (.DIODE(_1131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2890__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__A1 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A1 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__A1 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__A1 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2875__A1 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A1 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__A2 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__A2 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__A2 (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2859__A2 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2858__A2 (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__A (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2862__A2 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__A (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2863__A (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__A (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__A (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__A (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__A (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2864__A (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A0 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A0 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A0 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A0 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__A1 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3004__A1 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__A1 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__A1 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2877__A1 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2865__A1 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2870__B (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__A0 (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__A0 (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3019__A0 (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__A0 (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__A0 (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__A0 (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2925__A0 (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__A0 (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2901__A0 (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__A0 (.DIODE(_1239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__B (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__A (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__B (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__A (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2881__A (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__B (.DIODE(_1241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A (.DIODE(_1241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__A (.DIODE(_1241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__A (.DIODE(_1241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__A (.DIODE(_1241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__A (.DIODE(_1241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__A (.DIODE(_1241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__B (.DIODE(_1241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2924__A (.DIODE(_1241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__A (.DIODE(_1241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A (.DIODE(_1242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A (.DIODE(_1242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__B (.DIODE(_1242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__A (.DIODE(_1242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2934__B (.DIODE(_1242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2923__A (.DIODE(_1242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2912__A (.DIODE(_1242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2898__B (.DIODE(_1242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2883__D (.DIODE(_1242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__B (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__B (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3073__A0 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3064__A0 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3021__A0 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2969__A0 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2952__A0 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2938__A0 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__A0 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__A0 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2903__A0 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__A0 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__A0 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__A0 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3023__A0 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2971__A0 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__A0 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__A0 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2929__A0 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__A0 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__A0 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2891__A0 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3077__A0 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__A0 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__A0 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__A0 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A0 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__A0 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2931__A0 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2920__A0 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2907__A0 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2894__A0 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__A (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__A (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__B (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2897__A (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__B (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__B (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__B (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2900__A (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__A (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__B (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__A (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__B (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2900__B (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__A (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__A (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__B (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__C (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2913__A (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__B (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__B (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2935__A (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2912__B (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__B (.DIODE(_1271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__B (.DIODE(_1271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__A (.DIODE(_1271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A (.DIODE(_1271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__A (.DIODE(_1271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__A (.DIODE(_1271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3061__B (.DIODE(_1271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2924__B (.DIODE(_1271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__B (.DIODE(_1278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__B (.DIODE(_1278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(_1278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A (.DIODE(_1278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A (.DIODE(_1278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__A (.DIODE(_1278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__B (.DIODE(_1278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2935__B (.DIODE(_1278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__B (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B (.DIODE(_1287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A (.DIODE(_1287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__A (.DIODE(_1287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__B (.DIODE(_1287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__B (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__A (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__B (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__B (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__B (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2952__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__B (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__B (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__B (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__B (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__A (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__B (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__C (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__B (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__B (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__C (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__B (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__B (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__B (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__A (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__B (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3028__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A1 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__A1 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__A1 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A1 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__A1 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__A1 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3089__A1 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3080__A1 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__A1 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3033__A1 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__B (.DIODE(_1339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__B (.DIODE(_1339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A (.DIODE(_1339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__A (.DIODE(_1339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__B (.DIODE(_1339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__A1 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A1 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__A1 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A1 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__A1 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A1 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__A1 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A1 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__A (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__A (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3082__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3055__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__A1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__A1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__A (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3040__A (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__A1 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__A1 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__A1 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__A1 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__A1 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__A1 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3093__A1 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3084__A1 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__A1 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__A1 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__A1 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__A1 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__A1 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A1 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A1 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A1 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A1 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A1 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3332__A (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__A (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__B (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__A (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__B (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__B (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__A (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__B (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__B (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__B (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__A (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__A (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__B (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__B (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__B (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__B (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__B (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__B (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__S (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3093__S (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__S (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3089__S (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3200__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__A0 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__B (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__B (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__B (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__A (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__B (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__B (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__B (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__B (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__B (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__B (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__B (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__A0 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__A0 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__A0 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__A0 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__A0 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__A0 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__A0 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__A0 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__A0 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__A0 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__A0 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__A0 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A0 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3177__A0 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__A0 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__A0 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__A0 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3137__A0 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__A0 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__A0 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A0 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__A0 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A0 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3179__A0 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__A0 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3160__A0 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__A0 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__A0 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A0 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__A0 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__S (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__S (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__S (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__S (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__B (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__B (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__B (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__B (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__B (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__B (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__B (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__B (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__B (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__B (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__B (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__B (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__B (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__B (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__B (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__B (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__B (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__A (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__B (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__B (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__B (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__S (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__S (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__S (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__S (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3376__A0 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__A0 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__A0 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3316__A0 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__A0 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__A0 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__A0 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__A0 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__A0 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A0 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__A0 (.DIODE(_1458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__A0 (.DIODE(_1458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__A0 (.DIODE(_1458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__A0 (.DIODE(_1458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__A0 (.DIODE(_1458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__A0 (.DIODE(_1458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__A0 (.DIODE(_1458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__A0 (.DIODE(_1458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__A0 (.DIODE(_1458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A0 (.DIODE(_1458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__A0 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__A0 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__A0 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A0 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__A0 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__A0 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__A0 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__A0 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__A0 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__A0 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__B (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__B (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__B (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__B (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__B (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__B (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A1 (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A1 (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A1 (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__A1 (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__A1 (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__A1 (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A1 (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__A1 (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__A1 (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__A1 (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__A1 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A1 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__A1 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__A1 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__A1 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__A1 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__A1 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__A1 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3360__A1 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__A1 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3411__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3333__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__B (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__B (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__B (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__B (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__B (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__B (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__A (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__A0 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A0 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A0 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A0 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A0 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A0 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A0 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__A0 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A0 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__A0 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__A0 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__S (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__S (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__S (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__S (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A1 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A1 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A1 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A1 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A1 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__A1 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__A1 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A1 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A1 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A1 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__S (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__S (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__S (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__S (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A0 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A0 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A0 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A0 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A0 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A0 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A0 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__A0 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A0 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A0 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A0 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A0 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A0 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A0 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A0 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A0 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A0 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A0 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A0 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A0 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A0 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A0 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A0 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A0 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__A0 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A0 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A0 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A0 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__A0 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A0 (.DIODE(_1680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__B (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__S (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__S (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__S (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__S (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A1 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A1 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A1 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A1 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A1 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A1 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A1 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A1 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A1 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A1 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A0 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A0 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A0 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A0 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A0 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A0 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A0 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A0 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A0 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A0 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A0 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A0 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A0 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A0 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A0 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A0 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A0 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A0 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A0 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A0 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A0 (.DIODE(_1764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B (.DIODE(_1841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__D (.DIODE(_1841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__S (.DIODE(_1842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__S (.DIODE(_1842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__S (.DIODE(_1842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__S (.DIODE(_1842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__S (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__S (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__S (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__S (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__S (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__S (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__S (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__S (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__A0 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A0 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A0 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A0 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A0 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A0 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A0 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A0 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A0 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A0 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__A0 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A0 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__A0 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A0 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__A0 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A0 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A0 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A0 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A0 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A0 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__A0 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A0 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__A0 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A0 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__A0 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A0 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A0 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A0 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A0 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A0 (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A0 (.DIODE(_1874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A0 (.DIODE(_1874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__A0 (.DIODE(_1874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A0 (.DIODE(_1874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__A0 (.DIODE(_1874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A0 (.DIODE(_1874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A0 (.DIODE(_1874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A0 (.DIODE(_1874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__A0 (.DIODE(_1874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A0 (.DIODE(_1874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__S (.DIODE(_1896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__S (.DIODE(_1896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__S (.DIODE(_1896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__S (.DIODE(_1896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__B (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__C1 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__C1 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__C1 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__C1 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__C1 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__C1 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__C1 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__C1 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__C1 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__C1 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__A2 (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__A (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__A1 (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__A1 (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A1 (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__C (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A1 (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A_N (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__A0 (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__C1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__C1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__C1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__C1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__C1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__C1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__C1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__C1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__C1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__C1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__S (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__S (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__S (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__S (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__S (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__S (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__S (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__S (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__S (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__S (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__S (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__S (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A1 (.DIODE(chip_sel_override));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__A1 (.DIODE(chip_sel_override));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(oram_value[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(oram_value[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(oram_value[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(oram_value[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(oram_value[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(oram_value[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(oram_value[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(oram_value[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(oram_value[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(oram_value[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(oram_value[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(ram_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(ram_val[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(ram_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(ram_val[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(ram_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(ram_val[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(ram_val[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(ram_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(ram_val[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(ram_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(ram_val[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(ram_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(ram_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(ram_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(ram_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(ram_val[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(ram_val[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(ram_val[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(ram_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(ram_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(ram_val[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(ram_val[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(ram_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(ram_val[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(ram_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(ram_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(ram_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(ram_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(ram_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(ram_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(ram_val[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(ram_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A0 (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__A1 (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__B (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A_N (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__B (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A0 (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__B (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__A0 (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__A1 (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A1 (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__B (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A_N (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A0 (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__A (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__A0 (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__A3 (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A2 (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__B (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__B (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__A0 (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__B (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__D (.DIODE(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__A (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__A1 (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__B (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A1 (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A1 (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__B (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2543__D (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__B (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__B (.DIODE(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A1 (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__C (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2910__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2896__C (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__C_N (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__A_N (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__A1 (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A1 (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__C_N (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2910__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2896__A_N (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__A (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__A1 (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A1 (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__B (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__C (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__C (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__A_N (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2910__C_N (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2896__B (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__B (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__C (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2366__A1 (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__A (.DIODE(\tms1x00.wb_step ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__A (.DIODE(\tms1x00.wb_step ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__A1 (.DIODE(\tms1x00.wb_step ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__D (.DIODE(valid));
 sky130_fd_sc_hd__diode_2 ANTENNA__2368__B (.DIODE(valid));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__C (.DIODE(valid));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__C (.DIODE(valid));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__C (.DIODE(valid));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(wb_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(wbs_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(wbs_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(wbs_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(wbs_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(wbs_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(wbs_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(wbs_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(wbs_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(wbs_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(wbs_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(wbs_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(wbs_cyc_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(wbs_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(wbs_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(wbs_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(wbs_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(wbs_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(wbs_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(wbs_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(wbs_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(wbs_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(wbs_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2209__A0 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__A0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__A0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__A0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__2240__A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__2251__A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__2261__A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__2263__A0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__2265__A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__A0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__A0 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__2221__A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__2223__A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__2225__A0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__2227__A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__2208__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2291__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2293__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A_N (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__D_N (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2295__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__C (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__A_N (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__C_N (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2298__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2301__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__2303__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__2304__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2306__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2307__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2313__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2314__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__C (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__S (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2387__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__S (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__S (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__S (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__S (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__CLK (.DIODE(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__CLK (.DIODE(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_wb_clk_i_A (.DIODE(clknet_1_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_wb_clk_i_A (.DIODE(clknet_1_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_wb_clk_i_A (.DIODE(clknet_1_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_wb_clk_i_A (.DIODE(clknet_1_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_945 ();
 assign io_oeb[0] = net194;
 assign io_oeb[10] = net153;
 assign io_oeb[11] = net154;
 assign io_oeb[12] = net155;
 assign io_oeb[13] = net156;
 assign io_oeb[14] = net157;
 assign io_oeb[15] = net158;
 assign io_oeb[16] = net159;
 assign io_oeb[17] = net160;
 assign io_oeb[18] = net161;
 assign io_oeb[19] = net162;
 assign io_oeb[1] = net195;
 assign io_oeb[20] = net163;
 assign io_oeb[21] = net164;
 assign io_oeb[22] = net165;
 assign io_oeb[23] = net166;
 assign io_oeb[24] = net167;
 assign io_oeb[25] = net168;
 assign io_oeb[26] = net169;
 assign io_oeb[27] = net170;
 assign io_oeb[28] = net171;
 assign io_oeb[29] = net172;
 assign io_oeb[2] = net196;
 assign io_oeb[30] = net173;
 assign io_oeb[31] = net174;
 assign io_oeb[32] = net175;
 assign io_oeb[33] = net176;
 assign io_oeb[34] = net177;
 assign io_oeb[35] = net178;
 assign io_oeb[36] = net179;
 assign io_oeb[37] = net180;
 assign io_oeb[3] = net197;
 assign io_oeb[4] = net198;
 assign io_oeb[5] = net199;
 assign io_oeb[6] = net200;
 assign io_oeb[7] = net201;
 assign io_oeb[8] = net202;
 assign io_oeb[9] = net203;
 assign io_out[0] = net181;
 assign io_out[1] = net182;
 assign io_out[2] = net183;
 assign io_out[34] = net191;
 assign io_out[35] = net192;
 assign io_out[3] = net184;
 assign io_out[4] = net185;
 assign io_out[5] = net186;
 assign io_out[6] = net187;
 assign io_out[7] = net188;
 assign io_out[8] = net189;
 assign io_out[9] = net190;
 assign oram_addr[8] = net193;
endmodule

