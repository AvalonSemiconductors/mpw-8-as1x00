magic
tech sky130B
magscale 1 2
timestamp 1671146003
<< viali >>
rect 2789 6409 2823 6443
rect 1961 6273 1995 6307
rect 2605 6273 2639 6307
rect 3249 6273 3283 6307
rect 4445 6273 4479 6307
rect 5089 6273 5123 6307
rect 5733 6273 5767 6307
rect 9321 6273 9355 6307
rect 9781 6273 9815 6307
rect 3433 6137 3467 6171
rect 4629 6137 4663 6171
rect 2145 6069 2179 6103
rect 5273 6069 5307 6103
rect 9137 6069 9171 6103
rect 4813 5865 4847 5899
rect 3433 5797 3467 5831
rect 1869 5661 1903 5695
rect 2697 5661 2731 5695
rect 3249 5661 3283 5695
rect 4169 5661 4203 5695
rect 2053 5525 2087 5559
rect 2513 5525 2547 5559
rect 4353 5525 4387 5559
rect 2237 5321 2271 5355
rect 2881 5321 2915 5355
rect 3617 5321 3651 5355
rect 4169 5321 4203 5355
rect 1593 5185 1627 5219
rect 7205 5185 7239 5219
rect 1777 4981 1811 5015
rect 7389 4981 7423 5015
rect 1685 4777 1719 4811
rect 3157 4777 3191 4811
rect 2421 4573 2455 4607
rect 5549 4573 5583 4607
rect 7297 4573 7331 4607
rect 7941 4573 7975 4607
rect 2329 4437 2363 4471
rect 5733 4437 5767 4471
rect 7481 4437 7515 4471
rect 8125 4437 8159 4471
rect 1777 4097 1811 4131
rect 2697 4097 2731 4131
rect 4077 4097 4111 4131
rect 7481 4097 7515 4131
rect 7941 4097 7975 4131
rect 8585 4097 8619 4131
rect 2881 3893 2915 3927
rect 4261 3893 4295 3927
rect 7389 3893 7423 3927
rect 8125 3893 8159 3927
rect 8769 3893 8803 3927
rect 1593 3689 1627 3723
rect 7941 3485 7975 3519
rect 8125 3349 8159 3383
rect 14013 3009 14047 3043
rect 14197 2805 14231 2839
rect 1869 2397 1903 2431
rect 2513 2397 2547 2431
rect 3985 2397 4019 2431
rect 5273 2397 5307 2431
rect 6653 2397 6687 2431
rect 8033 2397 8067 2431
rect 9413 2397 9447 2431
rect 10793 2397 10827 2431
rect 12173 2397 12207 2431
rect 13461 2397 13495 2431
rect 1685 2261 1719 2295
rect 2697 2261 2731 2295
rect 4169 2261 4203 2295
rect 5457 2261 5491 2295
rect 6837 2261 6871 2295
rect 8217 2261 8251 2295
rect 9597 2261 9631 2295
rect 10977 2261 11011 2295
rect 12357 2261 12391 2295
rect 13645 2261 13679 2295
<< metal1 >>
rect 1104 6554 14971 6576
rect 1104 6502 4376 6554
rect 4428 6502 4440 6554
rect 4492 6502 4504 6554
rect 4556 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 7803 6554
rect 7855 6502 7867 6554
rect 7919 6502 7931 6554
rect 7983 6502 7995 6554
rect 8047 6502 8059 6554
rect 8111 6502 11230 6554
rect 11282 6502 11294 6554
rect 11346 6502 11358 6554
rect 11410 6502 11422 6554
rect 11474 6502 11486 6554
rect 11538 6502 14657 6554
rect 14709 6502 14721 6554
rect 14773 6502 14785 6554
rect 14837 6502 14849 6554
rect 14901 6502 14913 6554
rect 14965 6502 14971 6554
rect 1104 6480 14971 6502
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 6822 6440 6828 6452
rect 2823 6412 6828 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6304 2007 6307
rect 2222 6304 2228 6316
rect 1995 6276 2228 6304
rect 1995 6273 2007 6276
rect 1949 6267 2007 6273
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2498 6264 2504 6316
rect 2556 6304 2562 6316
rect 2593 6307 2651 6313
rect 2593 6304 2605 6307
rect 2556 6276 2605 6304
rect 2556 6264 2562 6276
rect 2593 6273 2605 6276
rect 2639 6304 2651 6307
rect 2682 6304 2688 6316
rect 2639 6276 2688 6304
rect 2639 6273 2651 6276
rect 2593 6267 2651 6273
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6304 3295 6307
rect 3602 6304 3608 6316
rect 3283 6276 3608 6304
rect 3283 6273 3295 6276
rect 3237 6267 3295 6273
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6304 4491 6307
rect 4706 6304 4712 6316
rect 4479 6276 4712 6304
rect 4479 6273 4491 6276
rect 4433 6267 4491 6273
rect 4706 6264 4712 6276
rect 4764 6264 4770 6316
rect 4982 6264 4988 6316
rect 5040 6304 5046 6316
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 5040 6276 5089 6304
rect 5040 6264 5046 6276
rect 5077 6273 5089 6276
rect 5123 6304 5135 6307
rect 5721 6307 5779 6313
rect 5721 6304 5733 6307
rect 5123 6276 5733 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 5721 6273 5733 6276
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 9309 6307 9367 6313
rect 9309 6304 9321 6307
rect 8720 6276 9321 6304
rect 8720 6264 8726 6276
rect 9309 6273 9321 6276
rect 9355 6304 9367 6307
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 9355 6276 9781 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 6638 6236 6644 6248
rect 3436 6208 6644 6236
rect 3436 6177 3464 6208
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 3421 6171 3479 6177
rect 3421 6137 3433 6171
rect 3467 6137 3479 6171
rect 3421 6131 3479 6137
rect 4617 6171 4675 6177
rect 4617 6137 4629 6171
rect 4663 6168 4675 6171
rect 6730 6168 6736 6180
rect 4663 6140 6736 6168
rect 4663 6137 4675 6140
rect 4617 6131 4675 6137
rect 6730 6128 6736 6140
rect 6788 6128 6794 6180
rect 2133 6103 2191 6109
rect 2133 6069 2145 6103
rect 2179 6100 2191 6103
rect 4062 6100 4068 6112
rect 2179 6072 4068 6100
rect 2179 6069 2191 6072
rect 2133 6063 2191 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 5261 6103 5319 6109
rect 5261 6069 5273 6103
rect 5307 6100 5319 6103
rect 5442 6100 5448 6112
rect 5307 6072 5448 6100
rect 5307 6069 5319 6072
rect 5261 6063 5319 6069
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 9125 6103 9183 6109
rect 9125 6100 9137 6103
rect 7616 6072 9137 6100
rect 7616 6060 7622 6072
rect 9125 6069 9137 6072
rect 9171 6069 9183 6103
rect 9125 6063 9183 6069
rect 1104 6010 14812 6032
rect 1104 5958 2663 6010
rect 2715 5958 2727 6010
rect 2779 5958 2791 6010
rect 2843 5958 2855 6010
rect 2907 5958 2919 6010
rect 2971 5958 6090 6010
rect 6142 5958 6154 6010
rect 6206 5958 6218 6010
rect 6270 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 9517 6010
rect 9569 5958 9581 6010
rect 9633 5958 9645 6010
rect 9697 5958 9709 6010
rect 9761 5958 9773 6010
rect 9825 5958 12944 6010
rect 12996 5958 13008 6010
rect 13060 5958 13072 6010
rect 13124 5958 13136 6010
rect 13188 5958 13200 6010
rect 13252 5958 14812 6010
rect 1104 5936 14812 5958
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 4801 5899 4859 5905
rect 4801 5896 4813 5899
rect 4764 5868 4813 5896
rect 4764 5856 4770 5868
rect 4801 5865 4813 5868
rect 4847 5865 4859 5899
rect 4801 5859 4859 5865
rect 3421 5831 3479 5837
rect 3421 5797 3433 5831
rect 3467 5828 3479 5831
rect 8570 5828 8576 5840
rect 3467 5800 8576 5828
rect 3467 5797 3479 5800
rect 3421 5791 3479 5797
rect 8570 5788 8576 5800
rect 8628 5788 8634 5840
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1820 5664 1869 5692
rect 1820 5652 1826 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2314 5652 2320 5704
rect 2372 5692 2378 5704
rect 2685 5695 2743 5701
rect 2685 5692 2697 5695
rect 2372 5664 2697 5692
rect 2372 5652 2378 5664
rect 2685 5661 2697 5664
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3237 5695 3295 5701
rect 3237 5692 3249 5695
rect 3200 5664 3249 5692
rect 3200 5652 3206 5664
rect 3237 5661 3249 5664
rect 3283 5661 3295 5695
rect 4154 5692 4160 5704
rect 4115 5664 4160 5692
rect 3237 5655 3295 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 2038 5556 2044 5568
rect 1999 5528 2044 5556
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 2406 5516 2412 5568
rect 2464 5556 2470 5568
rect 2501 5559 2559 5565
rect 2501 5556 2513 5559
rect 2464 5528 2513 5556
rect 2464 5516 2470 5528
rect 2501 5525 2513 5528
rect 2547 5525 2559 5559
rect 2501 5519 2559 5525
rect 4341 5559 4399 5565
rect 4341 5525 4353 5559
rect 4387 5556 4399 5559
rect 7650 5556 7656 5568
rect 4387 5528 7656 5556
rect 4387 5525 4399 5528
rect 4341 5519 4399 5525
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 1104 5466 14971 5488
rect 1104 5414 4376 5466
rect 4428 5414 4440 5466
rect 4492 5414 4504 5466
rect 4556 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 7803 5466
rect 7855 5414 7867 5466
rect 7919 5414 7931 5466
rect 7983 5414 7995 5466
rect 8047 5414 8059 5466
rect 8111 5414 11230 5466
rect 11282 5414 11294 5466
rect 11346 5414 11358 5466
rect 11410 5414 11422 5466
rect 11474 5414 11486 5466
rect 11538 5414 14657 5466
rect 14709 5414 14721 5466
rect 14773 5414 14785 5466
rect 14837 5414 14849 5466
rect 14901 5414 14913 5466
rect 14965 5414 14971 5466
rect 1104 5392 14971 5414
rect 2222 5352 2228 5364
rect 2183 5324 2228 5352
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 2869 5355 2927 5361
rect 2869 5352 2881 5355
rect 2556 5324 2881 5352
rect 2556 5312 2562 5324
rect 2869 5321 2881 5324
rect 2915 5321 2927 5355
rect 3602 5352 3608 5364
rect 3563 5324 3608 5352
rect 2869 5315 2927 5321
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 4154 5352 4160 5364
rect 4115 5324 4160 5352
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1578 5216 1584 5228
rect 1360 5188 1584 5216
rect 1360 5176 1366 5188
rect 1578 5176 1584 5188
rect 1636 5176 1642 5228
rect 6822 5176 6828 5228
rect 6880 5216 6886 5228
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 6880 5188 7205 5216
rect 6880 5176 6886 5188
rect 7193 5185 7205 5188
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 1765 5015 1823 5021
rect 1765 4981 1777 5015
rect 1811 5012 1823 5015
rect 2130 5012 2136 5024
rect 1811 4984 2136 5012
rect 1811 4981 1823 4984
rect 1765 4975 1823 4981
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 7374 5012 7380 5024
rect 7335 4984 7380 5012
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 1104 4922 14812 4944
rect 1104 4870 2663 4922
rect 2715 4870 2727 4922
rect 2779 4870 2791 4922
rect 2843 4870 2855 4922
rect 2907 4870 2919 4922
rect 2971 4870 6090 4922
rect 6142 4870 6154 4922
rect 6206 4870 6218 4922
rect 6270 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 9517 4922
rect 9569 4870 9581 4922
rect 9633 4870 9645 4922
rect 9697 4870 9709 4922
rect 9761 4870 9773 4922
rect 9825 4870 12944 4922
rect 12996 4870 13008 4922
rect 13060 4870 13072 4922
rect 13124 4870 13136 4922
rect 13188 4870 13200 4922
rect 13252 4870 14812 4922
rect 1104 4848 14812 4870
rect 842 4768 848 4820
rect 900 4808 906 4820
rect 1673 4811 1731 4817
rect 1673 4808 1685 4811
rect 900 4780 1685 4808
rect 900 4768 906 4780
rect 1673 4777 1685 4780
rect 1719 4808 1731 4811
rect 2314 4808 2320 4820
rect 1719 4780 2320 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 3142 4808 3148 4820
rect 3103 4780 3148 4808
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 6638 4632 6644 4684
rect 6696 4672 6702 4684
rect 6696 4644 7972 4672
rect 6696 4632 6702 4644
rect 2406 4604 2412 4616
rect 2367 4576 2412 4604
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 4062 4564 4068 4616
rect 4120 4604 4126 4616
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 4120 4576 5549 4604
rect 4120 4564 4126 4576
rect 5537 4573 5549 4576
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 7944 4613 7972 4644
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 6788 4576 7297 4604
rect 6788 4564 6794 4576
rect 7285 4573 7297 4576
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 2317 4471 2375 4477
rect 2317 4437 2329 4471
rect 2363 4468 2375 4471
rect 2498 4468 2504 4480
rect 2363 4440 2504 4468
rect 2363 4437 2375 4440
rect 2317 4431 2375 4437
rect 2498 4428 2504 4440
rect 2556 4428 2562 4480
rect 5721 4471 5779 4477
rect 5721 4437 5733 4471
rect 5767 4468 5779 4471
rect 6638 4468 6644 4480
rect 5767 4440 6644 4468
rect 5767 4437 5779 4440
rect 5721 4431 5779 4437
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 7466 4468 7472 4480
rect 7427 4440 7472 4468
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 8113 4471 8171 4477
rect 8113 4437 8125 4471
rect 8159 4468 8171 4471
rect 10778 4468 10784 4480
rect 8159 4440 10784 4468
rect 8159 4437 8171 4440
rect 8113 4431 8171 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 1104 4378 14971 4400
rect 1104 4326 4376 4378
rect 4428 4326 4440 4378
rect 4492 4326 4504 4378
rect 4556 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 7803 4378
rect 7855 4326 7867 4378
rect 7919 4326 7931 4378
rect 7983 4326 7995 4378
rect 8047 4326 8059 4378
rect 8111 4326 11230 4378
rect 11282 4326 11294 4378
rect 11346 4326 11358 4378
rect 11410 4326 11422 4378
rect 11474 4326 11486 4378
rect 11538 4326 14657 4378
rect 14709 4326 14721 4378
rect 14773 4326 14785 4378
rect 14837 4326 14849 4378
rect 14901 4326 14913 4378
rect 14965 4326 14971 4378
rect 1104 4304 14971 4326
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 13446 4264 13452 4276
rect 7524 4236 13452 4264
rect 7524 4224 7530 4236
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 1762 4128 1768 4140
rect 1723 4100 1768 4128
rect 1762 4088 1768 4100
rect 1820 4088 1826 4140
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2685 4131 2743 4137
rect 2685 4128 2697 4131
rect 2188 4100 2697 4128
rect 2188 4088 2194 4100
rect 2685 4097 2697 4100
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4097 4123 4131
rect 4065 4091 4123 4097
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 7558 4128 7564 4140
rect 7515 4100 7564 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 2038 4020 2044 4072
rect 2096 4060 2102 4072
rect 4080 4060 4108 4091
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 7650 4088 7656 4140
rect 7708 4128 7714 4140
rect 7929 4131 7987 4137
rect 7929 4128 7941 4131
rect 7708 4100 7941 4128
rect 7708 4088 7714 4100
rect 7929 4097 7941 4100
rect 7975 4097 7987 4131
rect 8570 4128 8576 4140
rect 8531 4100 8576 4128
rect 7929 4091 7987 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 2096 4032 4108 4060
rect 2096 4020 2102 4032
rect 2869 3927 2927 3933
rect 2869 3893 2881 3927
rect 2915 3924 2927 3927
rect 3970 3924 3976 3936
rect 2915 3896 3976 3924
rect 2915 3893 2927 3896
rect 2869 3887 2927 3893
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3924 4307 3927
rect 5258 3924 5264 3936
rect 4295 3896 5264 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7377 3927 7435 3933
rect 7377 3924 7389 3927
rect 6972 3896 7389 3924
rect 6972 3884 6978 3896
rect 7377 3893 7389 3896
rect 7423 3893 7435 3927
rect 7377 3887 7435 3893
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8662 3924 8668 3936
rect 8159 3896 8668 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 8757 3927 8815 3933
rect 8757 3893 8769 3927
rect 8803 3924 8815 3927
rect 9398 3924 9404 3936
rect 8803 3896 9404 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 1104 3834 14812 3856
rect 1104 3782 2663 3834
rect 2715 3782 2727 3834
rect 2779 3782 2791 3834
rect 2843 3782 2855 3834
rect 2907 3782 2919 3834
rect 2971 3782 6090 3834
rect 6142 3782 6154 3834
rect 6206 3782 6218 3834
rect 6270 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 9517 3834
rect 9569 3782 9581 3834
rect 9633 3782 9645 3834
rect 9697 3782 9709 3834
rect 9761 3782 9773 3834
rect 9825 3782 12944 3834
rect 12996 3782 13008 3834
rect 13060 3782 13072 3834
rect 13124 3782 13136 3834
rect 13188 3782 13200 3834
rect 13252 3782 14812 3834
rect 1104 3760 14812 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 5500 3488 7941 3516
rect 5500 3476 5506 3488
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 8113 3383 8171 3389
rect 8113 3349 8125 3383
rect 8159 3380 8171 3383
rect 13998 3380 14004 3392
rect 8159 3352 14004 3380
rect 8159 3349 8171 3352
rect 8113 3343 8171 3349
rect 13998 3340 14004 3352
rect 14056 3340 14062 3392
rect 1104 3290 14971 3312
rect 1104 3238 4376 3290
rect 4428 3238 4440 3290
rect 4492 3238 4504 3290
rect 4556 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 7803 3290
rect 7855 3238 7867 3290
rect 7919 3238 7931 3290
rect 7983 3238 7995 3290
rect 8047 3238 8059 3290
rect 8111 3238 11230 3290
rect 11282 3238 11294 3290
rect 11346 3238 11358 3290
rect 11410 3238 11422 3290
rect 11474 3238 11486 3290
rect 11538 3238 14657 3290
rect 14709 3238 14721 3290
rect 14773 3238 14785 3290
rect 14837 3238 14849 3290
rect 14901 3238 14913 3290
rect 14965 3238 14971 3290
rect 1104 3216 14971 3238
rect 13998 3040 14004 3052
rect 13959 3012 14004 3040
rect 13998 3000 14004 3012
rect 14056 3000 14062 3052
rect 14185 2839 14243 2845
rect 14185 2805 14197 2839
rect 14231 2836 14243 2839
rect 14550 2836 14556 2848
rect 14231 2808 14556 2836
rect 14231 2805 14243 2808
rect 14185 2799 14243 2805
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 1104 2746 14812 2768
rect 1104 2694 2663 2746
rect 2715 2694 2727 2746
rect 2779 2694 2791 2746
rect 2843 2694 2855 2746
rect 2907 2694 2919 2746
rect 2971 2694 6090 2746
rect 6142 2694 6154 2746
rect 6206 2694 6218 2746
rect 6270 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 9517 2746
rect 9569 2694 9581 2746
rect 9633 2694 9645 2746
rect 9697 2694 9709 2746
rect 9761 2694 9773 2746
rect 9825 2694 12944 2746
rect 12996 2694 13008 2746
rect 13060 2694 13072 2746
rect 13124 2694 13136 2746
rect 13188 2694 13200 2746
rect 13252 2694 14812 2746
rect 1104 2672 14812 2694
rect 6914 2496 6920 2508
rect 1872 2468 6920 2496
rect 1872 2437 1900 2468
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 8662 2456 8668 2508
rect 8720 2496 8726 2508
rect 8720 2468 12204 2496
rect 8720 2456 8726 2468
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 2498 2428 2504 2440
rect 2459 2400 2504 2428
rect 1857 2391 1915 2397
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 3970 2428 3976 2440
rect 3931 2400 3976 2428
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 5258 2428 5264 2440
rect 5219 2400 5264 2428
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 6638 2428 6644 2440
rect 6599 2400 6644 2428
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 7374 2388 7380 2440
rect 7432 2428 7438 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7432 2400 8033 2428
rect 7432 2388 7438 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 9398 2428 9404 2440
rect 9359 2400 9404 2428
rect 8021 2391 8079 2397
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 10778 2428 10784 2440
rect 10739 2400 10784 2428
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 12176 2437 12204 2468
rect 12161 2431 12219 2437
rect 12161 2397 12173 2431
rect 12207 2397 12219 2431
rect 13446 2428 13452 2440
rect 13407 2400 13452 2428
rect 12161 2391 12219 2397
rect 13446 2388 13452 2400
rect 13504 2388 13510 2440
rect 1026 2252 1032 2304
rect 1084 2292 1090 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1084 2264 1685 2292
rect 1084 2252 1090 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 2406 2252 2412 2304
rect 2464 2292 2470 2304
rect 2685 2295 2743 2301
rect 2685 2292 2697 2295
rect 2464 2264 2697 2292
rect 2464 2252 2470 2264
rect 2685 2261 2697 2264
rect 2731 2261 2743 2295
rect 2685 2255 2743 2261
rect 3786 2252 3792 2304
rect 3844 2292 3850 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 3844 2264 4169 2292
rect 3844 2252 3850 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5224 2264 5457 2292
rect 5224 2252 5230 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 6546 2252 6552 2304
rect 6604 2292 6610 2304
rect 6825 2295 6883 2301
rect 6825 2292 6837 2295
rect 6604 2264 6837 2292
rect 6604 2252 6610 2264
rect 6825 2261 6837 2264
rect 6871 2261 6883 2295
rect 8202 2292 8208 2304
rect 8163 2264 8208 2292
rect 6825 2255 6883 2261
rect 8202 2252 8208 2264
rect 8260 2252 8266 2304
rect 9306 2252 9312 2304
rect 9364 2292 9370 2304
rect 9585 2295 9643 2301
rect 9585 2292 9597 2295
rect 9364 2264 9597 2292
rect 9364 2252 9370 2264
rect 9585 2261 9597 2264
rect 9631 2261 9643 2295
rect 9585 2255 9643 2261
rect 10686 2252 10692 2304
rect 10744 2292 10750 2304
rect 10965 2295 11023 2301
rect 10965 2292 10977 2295
rect 10744 2264 10977 2292
rect 10744 2252 10750 2264
rect 10965 2261 10977 2264
rect 11011 2261 11023 2295
rect 10965 2255 11023 2261
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 12345 2295 12403 2301
rect 12345 2292 12357 2295
rect 12124 2264 12357 2292
rect 12124 2252 12130 2264
rect 12345 2261 12357 2264
rect 12391 2261 12403 2295
rect 12345 2255 12403 2261
rect 13446 2252 13452 2304
rect 13504 2292 13510 2304
rect 13633 2295 13691 2301
rect 13633 2292 13645 2295
rect 13504 2264 13645 2292
rect 13504 2252 13510 2264
rect 13633 2261 13645 2264
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 1104 2202 14971 2224
rect 1104 2150 4376 2202
rect 4428 2150 4440 2202
rect 4492 2150 4504 2202
rect 4556 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 7803 2202
rect 7855 2150 7867 2202
rect 7919 2150 7931 2202
rect 7983 2150 7995 2202
rect 8047 2150 8059 2202
rect 8111 2150 11230 2202
rect 11282 2150 11294 2202
rect 11346 2150 11358 2202
rect 11410 2150 11422 2202
rect 11474 2150 11486 2202
rect 11538 2150 14657 2202
rect 14709 2150 14721 2202
rect 14773 2150 14785 2202
rect 14837 2150 14849 2202
rect 14901 2150 14913 2202
rect 14965 2150 14971 2202
rect 1104 2128 14971 2150
<< via1 >>
rect 4376 6502 4428 6554
rect 4440 6502 4492 6554
rect 4504 6502 4556 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 7803 6502 7855 6554
rect 7867 6502 7919 6554
rect 7931 6502 7983 6554
rect 7995 6502 8047 6554
rect 8059 6502 8111 6554
rect 11230 6502 11282 6554
rect 11294 6502 11346 6554
rect 11358 6502 11410 6554
rect 11422 6502 11474 6554
rect 11486 6502 11538 6554
rect 14657 6502 14709 6554
rect 14721 6502 14773 6554
rect 14785 6502 14837 6554
rect 14849 6502 14901 6554
rect 14913 6502 14965 6554
rect 6828 6400 6880 6452
rect 2228 6264 2280 6316
rect 2504 6264 2556 6316
rect 2688 6264 2740 6316
rect 3608 6264 3660 6316
rect 4712 6264 4764 6316
rect 4988 6264 5040 6316
rect 8668 6264 8720 6316
rect 6644 6196 6696 6248
rect 6736 6128 6788 6180
rect 4068 6060 4120 6112
rect 5448 6060 5500 6112
rect 7564 6060 7616 6112
rect 2663 5958 2715 6010
rect 2727 5958 2779 6010
rect 2791 5958 2843 6010
rect 2855 5958 2907 6010
rect 2919 5958 2971 6010
rect 6090 5958 6142 6010
rect 6154 5958 6206 6010
rect 6218 5958 6270 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 9517 5958 9569 6010
rect 9581 5958 9633 6010
rect 9645 5958 9697 6010
rect 9709 5958 9761 6010
rect 9773 5958 9825 6010
rect 12944 5958 12996 6010
rect 13008 5958 13060 6010
rect 13072 5958 13124 6010
rect 13136 5958 13188 6010
rect 13200 5958 13252 6010
rect 4712 5856 4764 5908
rect 8576 5788 8628 5840
rect 1768 5652 1820 5704
rect 2320 5652 2372 5704
rect 3148 5652 3200 5704
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 2044 5559 2096 5568
rect 2044 5525 2053 5559
rect 2053 5525 2087 5559
rect 2087 5525 2096 5559
rect 2044 5516 2096 5525
rect 2412 5516 2464 5568
rect 7656 5516 7708 5568
rect 4376 5414 4428 5466
rect 4440 5414 4492 5466
rect 4504 5414 4556 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 7803 5414 7855 5466
rect 7867 5414 7919 5466
rect 7931 5414 7983 5466
rect 7995 5414 8047 5466
rect 8059 5414 8111 5466
rect 11230 5414 11282 5466
rect 11294 5414 11346 5466
rect 11358 5414 11410 5466
rect 11422 5414 11474 5466
rect 11486 5414 11538 5466
rect 14657 5414 14709 5466
rect 14721 5414 14773 5466
rect 14785 5414 14837 5466
rect 14849 5414 14901 5466
rect 14913 5414 14965 5466
rect 2228 5355 2280 5364
rect 2228 5321 2237 5355
rect 2237 5321 2271 5355
rect 2271 5321 2280 5355
rect 2228 5312 2280 5321
rect 2504 5312 2556 5364
rect 3608 5355 3660 5364
rect 3608 5321 3617 5355
rect 3617 5321 3651 5355
rect 3651 5321 3660 5355
rect 3608 5312 3660 5321
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4160 5312 4212 5321
rect 1308 5176 1360 5228
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 6828 5176 6880 5228
rect 2136 4972 2188 5024
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 2663 4870 2715 4922
rect 2727 4870 2779 4922
rect 2791 4870 2843 4922
rect 2855 4870 2907 4922
rect 2919 4870 2971 4922
rect 6090 4870 6142 4922
rect 6154 4870 6206 4922
rect 6218 4870 6270 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 9517 4870 9569 4922
rect 9581 4870 9633 4922
rect 9645 4870 9697 4922
rect 9709 4870 9761 4922
rect 9773 4870 9825 4922
rect 12944 4870 12996 4922
rect 13008 4870 13060 4922
rect 13072 4870 13124 4922
rect 13136 4870 13188 4922
rect 13200 4870 13252 4922
rect 848 4768 900 4820
rect 2320 4768 2372 4820
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 6644 4632 6696 4684
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 4068 4564 4120 4616
rect 6736 4564 6788 4616
rect 2504 4428 2556 4480
rect 6644 4428 6696 4480
rect 7472 4471 7524 4480
rect 7472 4437 7481 4471
rect 7481 4437 7515 4471
rect 7515 4437 7524 4471
rect 7472 4428 7524 4437
rect 10784 4428 10836 4480
rect 4376 4326 4428 4378
rect 4440 4326 4492 4378
rect 4504 4326 4556 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 7803 4326 7855 4378
rect 7867 4326 7919 4378
rect 7931 4326 7983 4378
rect 7995 4326 8047 4378
rect 8059 4326 8111 4378
rect 11230 4326 11282 4378
rect 11294 4326 11346 4378
rect 11358 4326 11410 4378
rect 11422 4326 11474 4378
rect 11486 4326 11538 4378
rect 14657 4326 14709 4378
rect 14721 4326 14773 4378
rect 14785 4326 14837 4378
rect 14849 4326 14901 4378
rect 14913 4326 14965 4378
rect 7472 4224 7524 4276
rect 13452 4224 13504 4276
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 2136 4088 2188 4140
rect 2044 4020 2096 4072
rect 7564 4088 7616 4140
rect 7656 4088 7708 4140
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 3976 3884 4028 3936
rect 5264 3884 5316 3936
rect 6920 3884 6972 3936
rect 8668 3884 8720 3936
rect 9404 3884 9456 3936
rect 2663 3782 2715 3834
rect 2727 3782 2779 3834
rect 2791 3782 2843 3834
rect 2855 3782 2907 3834
rect 2919 3782 2971 3834
rect 6090 3782 6142 3834
rect 6154 3782 6206 3834
rect 6218 3782 6270 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 9517 3782 9569 3834
rect 9581 3782 9633 3834
rect 9645 3782 9697 3834
rect 9709 3782 9761 3834
rect 9773 3782 9825 3834
rect 12944 3782 12996 3834
rect 13008 3782 13060 3834
rect 13072 3782 13124 3834
rect 13136 3782 13188 3834
rect 13200 3782 13252 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 5448 3476 5500 3528
rect 14004 3340 14056 3392
rect 4376 3238 4428 3290
rect 4440 3238 4492 3290
rect 4504 3238 4556 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 7803 3238 7855 3290
rect 7867 3238 7919 3290
rect 7931 3238 7983 3290
rect 7995 3238 8047 3290
rect 8059 3238 8111 3290
rect 11230 3238 11282 3290
rect 11294 3238 11346 3290
rect 11358 3238 11410 3290
rect 11422 3238 11474 3290
rect 11486 3238 11538 3290
rect 14657 3238 14709 3290
rect 14721 3238 14773 3290
rect 14785 3238 14837 3290
rect 14849 3238 14901 3290
rect 14913 3238 14965 3290
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 14556 2796 14608 2848
rect 2663 2694 2715 2746
rect 2727 2694 2779 2746
rect 2791 2694 2843 2746
rect 2855 2694 2907 2746
rect 2919 2694 2971 2746
rect 6090 2694 6142 2746
rect 6154 2694 6206 2746
rect 6218 2694 6270 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 9517 2694 9569 2746
rect 9581 2694 9633 2746
rect 9645 2694 9697 2746
rect 9709 2694 9761 2746
rect 9773 2694 9825 2746
rect 12944 2694 12996 2746
rect 13008 2694 13060 2746
rect 13072 2694 13124 2746
rect 13136 2694 13188 2746
rect 13200 2694 13252 2746
rect 6920 2456 6972 2508
rect 8668 2456 8720 2508
rect 2504 2431 2556 2440
rect 2504 2397 2513 2431
rect 2513 2397 2547 2431
rect 2547 2397 2556 2431
rect 2504 2388 2556 2397
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 7380 2388 7432 2440
rect 9404 2431 9456 2440
rect 9404 2397 9413 2431
rect 9413 2397 9447 2431
rect 9447 2397 9456 2431
rect 9404 2388 9456 2397
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 13452 2431 13504 2440
rect 13452 2397 13461 2431
rect 13461 2397 13495 2431
rect 13495 2397 13504 2431
rect 13452 2388 13504 2397
rect 1032 2252 1084 2304
rect 2412 2252 2464 2304
rect 3792 2252 3844 2304
rect 5172 2252 5224 2304
rect 6552 2252 6604 2304
rect 8208 2295 8260 2304
rect 8208 2261 8217 2295
rect 8217 2261 8251 2295
rect 8251 2261 8260 2295
rect 8208 2252 8260 2261
rect 9312 2252 9364 2304
rect 10692 2252 10744 2304
rect 12072 2252 12124 2304
rect 13452 2252 13504 2304
rect 4376 2150 4428 2202
rect 4440 2150 4492 2202
rect 4504 2150 4556 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 7803 2150 7855 2202
rect 7867 2150 7919 2202
rect 7931 2150 7983 2202
rect 7995 2150 8047 2202
rect 8059 2150 8111 2202
rect 11230 2150 11282 2202
rect 11294 2150 11346 2202
rect 11358 2150 11410 2202
rect 11422 2150 11474 2202
rect 11486 2150 11538 2202
rect 14657 2150 14709 2202
rect 14721 2150 14773 2202
rect 14785 2150 14837 2202
rect 14849 2150 14901 2202
rect 14913 2150 14965 2202
<< metal2 >>
rect 386 8200 442 9000
rect 846 8200 902 9000
rect 1306 8200 1362 9000
rect 1766 8200 1822 9000
rect 2226 8200 2282 9000
rect 2686 8200 2742 9000
rect 3146 8200 3202 9000
rect 3606 8200 3662 9000
rect 4066 8200 4122 9000
rect 4526 8200 4582 9000
rect 4986 8200 5042 9000
rect 5446 8200 5502 9000
rect 5906 8200 5962 9000
rect 6366 8200 6422 9000
rect 6826 8200 6882 9000
rect 7286 8200 7342 9000
rect 7746 8200 7802 9000
rect 8206 8200 8262 9000
rect 8666 8200 8722 9000
rect 9126 8200 9182 9000
rect 9586 8200 9642 9000
rect 10046 8200 10102 9000
rect 10506 8200 10562 9000
rect 10966 8200 11022 9000
rect 11426 8200 11482 9000
rect 11886 8200 11942 9000
rect 12346 8200 12402 9000
rect 12806 8200 12862 9000
rect 13266 8200 13322 9000
rect 13726 8200 13782 9000
rect 14186 8200 14242 9000
rect 14646 8200 14702 9000
rect 15106 8200 15162 9000
rect 15566 8200 15622 9000
rect 860 4826 888 8200
rect 1320 5234 1348 8200
rect 1780 5710 1808 8200
rect 2240 6322 2268 8200
rect 2700 6322 2728 8200
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 848 4820 900 4826
rect 848 4762 900 4768
rect 1596 3738 1624 5170
rect 1780 4146 1808 5646
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 2056 4078 2084 5510
rect 2240 5370 2268 6258
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2148 4146 2176 4966
rect 2332 4826 2360 5646
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2424 4622 2452 5510
rect 2516 5370 2544 6258
rect 2663 6012 2971 6021
rect 2663 6010 2669 6012
rect 2725 6010 2749 6012
rect 2805 6010 2829 6012
rect 2885 6010 2909 6012
rect 2965 6010 2971 6012
rect 2725 5958 2727 6010
rect 2907 5958 2909 6010
rect 2663 5956 2669 5958
rect 2725 5956 2749 5958
rect 2805 5956 2829 5958
rect 2885 5956 2909 5958
rect 2965 5956 2971 5958
rect 2663 5947 2971 5956
rect 3160 5710 3188 8200
rect 3620 6322 3648 8200
rect 4080 6338 4108 8200
rect 4540 6746 4568 8200
rect 4540 6718 4752 6746
rect 4376 6556 4684 6565
rect 4376 6554 4382 6556
rect 4438 6554 4462 6556
rect 4518 6554 4542 6556
rect 4598 6554 4622 6556
rect 4678 6554 4684 6556
rect 4438 6502 4440 6554
rect 4620 6502 4622 6554
rect 4376 6500 4382 6502
rect 4438 6500 4462 6502
rect 4518 6500 4542 6502
rect 4598 6500 4622 6502
rect 4678 6500 4684 6502
rect 4376 6491 4684 6500
rect 3608 6316 3660 6322
rect 4080 6310 4200 6338
rect 4724 6322 4752 6718
rect 5000 6322 5028 8200
rect 7803 6556 8111 6565
rect 7803 6554 7809 6556
rect 7865 6554 7889 6556
rect 7945 6554 7969 6556
rect 8025 6554 8049 6556
rect 8105 6554 8111 6556
rect 7865 6502 7867 6554
rect 8047 6502 8049 6554
rect 7803 6500 7809 6502
rect 7865 6500 7889 6502
rect 7945 6500 7969 6502
rect 8025 6500 8049 6502
rect 8105 6500 8111 6502
rect 7803 6491 8111 6500
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 3608 6258 3660 6264
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2663 4924 2971 4933
rect 2663 4922 2669 4924
rect 2725 4922 2749 4924
rect 2805 4922 2829 4924
rect 2885 4922 2909 4924
rect 2965 4922 2971 4924
rect 2725 4870 2727 4922
rect 2907 4870 2909 4922
rect 2663 4868 2669 4870
rect 2725 4868 2749 4870
rect 2805 4868 2829 4870
rect 2885 4868 2909 4870
rect 2965 4868 2971 4870
rect 2663 4859 2971 4868
rect 3160 4826 3188 5646
rect 3620 5370 3648 6258
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 4080 4622 4108 6054
rect 4172 5710 4200 6310
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 4724 5914 4752 6258
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4172 5370 4200 5646
rect 4376 5468 4684 5477
rect 4376 5466 4382 5468
rect 4438 5466 4462 5468
rect 4518 5466 4542 5468
rect 4598 5466 4622 5468
rect 4678 5466 4684 5468
rect 4438 5414 4440 5466
rect 4620 5414 4622 5466
rect 4376 5412 4382 5414
rect 4438 5412 4462 5414
rect 4518 5412 4542 5414
rect 4598 5412 4622 5414
rect 4678 5412 4684 5414
rect 4376 5403 4684 5412
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 2516 2446 2544 4422
rect 4376 4380 4684 4389
rect 4376 4378 4382 4380
rect 4438 4378 4462 4380
rect 4518 4378 4542 4380
rect 4598 4378 4622 4380
rect 4678 4378 4684 4380
rect 4438 4326 4440 4378
rect 4620 4326 4622 4378
rect 4376 4324 4382 4326
rect 4438 4324 4462 4326
rect 4518 4324 4542 4326
rect 4598 4324 4622 4326
rect 4678 4324 4684 4326
rect 4376 4315 4684 4324
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 2663 3836 2971 3845
rect 2663 3834 2669 3836
rect 2725 3834 2749 3836
rect 2805 3834 2829 3836
rect 2885 3834 2909 3836
rect 2965 3834 2971 3836
rect 2725 3782 2727 3834
rect 2907 3782 2909 3834
rect 2663 3780 2669 3782
rect 2725 3780 2749 3782
rect 2805 3780 2829 3782
rect 2885 3780 2909 3782
rect 2965 3780 2971 3782
rect 2663 3771 2971 3780
rect 2663 2748 2971 2757
rect 2663 2746 2669 2748
rect 2725 2746 2749 2748
rect 2805 2746 2829 2748
rect 2885 2746 2909 2748
rect 2965 2746 2971 2748
rect 2725 2694 2727 2746
rect 2907 2694 2909 2746
rect 2663 2692 2669 2694
rect 2725 2692 2749 2694
rect 2805 2692 2829 2694
rect 2885 2692 2909 2694
rect 2965 2692 2971 2694
rect 2663 2683 2971 2692
rect 3988 2446 4016 3878
rect 4376 3292 4684 3301
rect 4376 3290 4382 3292
rect 4438 3290 4462 3292
rect 4518 3290 4542 3292
rect 4598 3290 4622 3292
rect 4678 3290 4684 3292
rect 4438 3238 4440 3290
rect 4620 3238 4622 3290
rect 4376 3236 4382 3238
rect 4438 3236 4462 3238
rect 4518 3236 4542 3238
rect 4598 3236 4622 3238
rect 4678 3236 4684 3238
rect 4376 3227 4684 3236
rect 5276 2446 5304 3878
rect 5460 3534 5488 6054
rect 6090 6012 6398 6021
rect 6090 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6336 6012
rect 6392 6010 6398 6012
rect 6152 5958 6154 6010
rect 6334 5958 6336 6010
rect 6090 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6336 5958
rect 6392 5956 6398 5958
rect 6090 5947 6398 5956
rect 6090 4924 6398 4933
rect 6090 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6336 4924
rect 6392 4922 6398 4924
rect 6152 4870 6154 4922
rect 6334 4870 6336 4922
rect 6090 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6336 4870
rect 6392 4868 6398 4870
rect 6090 4859 6398 4868
rect 6656 4690 6684 6190
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6748 4622 6776 6122
rect 6840 5234 6868 6394
rect 8680 6322 8708 8200
rect 11230 6556 11538 6565
rect 11230 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11396 6556
rect 11452 6554 11476 6556
rect 11532 6554 11538 6556
rect 11292 6502 11294 6554
rect 11474 6502 11476 6554
rect 11230 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11396 6502
rect 11452 6500 11476 6502
rect 11532 6500 11538 6502
rect 11230 6491 11538 6500
rect 14657 6556 14965 6565
rect 14657 6554 14663 6556
rect 14719 6554 14743 6556
rect 14799 6554 14823 6556
rect 14879 6554 14903 6556
rect 14959 6554 14965 6556
rect 14719 6502 14721 6554
rect 14901 6502 14903 6554
rect 14657 6500 14663 6502
rect 14719 6500 14743 6502
rect 14799 6500 14823 6502
rect 14879 6500 14903 6502
rect 14959 6500 14965 6502
rect 14657 6491 14965 6500
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6090 3836 6398 3845
rect 6090 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6336 3836
rect 6392 3834 6398 3836
rect 6152 3782 6154 3834
rect 6334 3782 6336 3834
rect 6090 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6336 3782
rect 6392 3780 6398 3782
rect 6090 3771 6398 3780
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 6090 2748 6398 2757
rect 6090 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6336 2748
rect 6392 2746 6398 2748
rect 6152 2694 6154 2746
rect 6334 2694 6336 2746
rect 6090 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6336 2694
rect 6392 2692 6398 2694
rect 6090 2683 6398 2692
rect 6656 2446 6684 4422
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6932 2514 6960 3878
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7392 2446 7420 4966
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7484 4282 7512 4422
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7576 4146 7604 6054
rect 9517 6012 9825 6021
rect 9517 6010 9523 6012
rect 9579 6010 9603 6012
rect 9659 6010 9683 6012
rect 9739 6010 9763 6012
rect 9819 6010 9825 6012
rect 9579 5958 9581 6010
rect 9761 5958 9763 6010
rect 9517 5956 9523 5958
rect 9579 5956 9603 5958
rect 9659 5956 9683 5958
rect 9739 5956 9763 5958
rect 9819 5956 9825 5958
rect 9517 5947 9825 5956
rect 12944 6012 13252 6021
rect 12944 6010 12950 6012
rect 13006 6010 13030 6012
rect 13086 6010 13110 6012
rect 13166 6010 13190 6012
rect 13246 6010 13252 6012
rect 13006 5958 13008 6010
rect 13188 5958 13190 6010
rect 12944 5956 12950 5958
rect 13006 5956 13030 5958
rect 13086 5956 13110 5958
rect 13166 5956 13190 5958
rect 13246 5956 13252 5958
rect 12944 5947 13252 5956
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7668 4146 7696 5510
rect 7803 5468 8111 5477
rect 7803 5466 7809 5468
rect 7865 5466 7889 5468
rect 7945 5466 7969 5468
rect 8025 5466 8049 5468
rect 8105 5466 8111 5468
rect 7865 5414 7867 5466
rect 8047 5414 8049 5466
rect 7803 5412 7809 5414
rect 7865 5412 7889 5414
rect 7945 5412 7969 5414
rect 8025 5412 8049 5414
rect 8105 5412 8111 5414
rect 7803 5403 8111 5412
rect 7803 4380 8111 4389
rect 7803 4378 7809 4380
rect 7865 4378 7889 4380
rect 7945 4378 7969 4380
rect 8025 4378 8049 4380
rect 8105 4378 8111 4380
rect 7865 4326 7867 4378
rect 8047 4326 8049 4378
rect 7803 4324 7809 4326
rect 7865 4324 7889 4326
rect 7945 4324 7969 4326
rect 8025 4324 8049 4326
rect 8105 4324 8111 4326
rect 7803 4315 8111 4324
rect 8588 4146 8616 5782
rect 11230 5468 11538 5477
rect 11230 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11396 5468
rect 11452 5466 11476 5468
rect 11532 5466 11538 5468
rect 11292 5414 11294 5466
rect 11474 5414 11476 5466
rect 11230 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11396 5414
rect 11452 5412 11476 5414
rect 11532 5412 11538 5414
rect 11230 5403 11538 5412
rect 14657 5468 14965 5477
rect 14657 5466 14663 5468
rect 14719 5466 14743 5468
rect 14799 5466 14823 5468
rect 14879 5466 14903 5468
rect 14959 5466 14965 5468
rect 14719 5414 14721 5466
rect 14901 5414 14903 5466
rect 14657 5412 14663 5414
rect 14719 5412 14743 5414
rect 14799 5412 14823 5414
rect 14879 5412 14903 5414
rect 14959 5412 14965 5414
rect 14657 5403 14965 5412
rect 9517 4924 9825 4933
rect 9517 4922 9523 4924
rect 9579 4922 9603 4924
rect 9659 4922 9683 4924
rect 9739 4922 9763 4924
rect 9819 4922 9825 4924
rect 9579 4870 9581 4922
rect 9761 4870 9763 4922
rect 9517 4868 9523 4870
rect 9579 4868 9603 4870
rect 9659 4868 9683 4870
rect 9739 4868 9763 4870
rect 9819 4868 9825 4870
rect 9517 4859 9825 4868
rect 12944 4924 13252 4933
rect 12944 4922 12950 4924
rect 13006 4922 13030 4924
rect 13086 4922 13110 4924
rect 13166 4922 13190 4924
rect 13246 4922 13252 4924
rect 13006 4870 13008 4922
rect 13188 4870 13190 4922
rect 12944 4868 12950 4870
rect 13006 4868 13030 4870
rect 13086 4868 13110 4870
rect 13166 4868 13190 4870
rect 13246 4868 13252 4870
rect 12944 4859 13252 4868
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 7803 3292 8111 3301
rect 7803 3290 7809 3292
rect 7865 3290 7889 3292
rect 7945 3290 7969 3292
rect 8025 3290 8049 3292
rect 8105 3290 8111 3292
rect 7865 3238 7867 3290
rect 8047 3238 8049 3290
rect 7803 3236 7809 3238
rect 7865 3236 7889 3238
rect 7945 3236 7969 3238
rect 8025 3236 8049 3238
rect 8105 3236 8111 3238
rect 7803 3227 8111 3236
rect 8680 2514 8708 3878
rect 8668 2508 8720 2514
rect 8668 2450 8720 2456
rect 9416 2446 9444 3878
rect 9517 3836 9825 3845
rect 9517 3834 9523 3836
rect 9579 3834 9603 3836
rect 9659 3834 9683 3836
rect 9739 3834 9763 3836
rect 9819 3834 9825 3836
rect 9579 3782 9581 3834
rect 9761 3782 9763 3834
rect 9517 3780 9523 3782
rect 9579 3780 9603 3782
rect 9659 3780 9683 3782
rect 9739 3780 9763 3782
rect 9819 3780 9825 3782
rect 9517 3771 9825 3780
rect 9517 2748 9825 2757
rect 9517 2746 9523 2748
rect 9579 2746 9603 2748
rect 9659 2746 9683 2748
rect 9739 2746 9763 2748
rect 9819 2746 9825 2748
rect 9579 2694 9581 2746
rect 9761 2694 9763 2746
rect 9517 2692 9523 2694
rect 9579 2692 9603 2694
rect 9659 2692 9683 2694
rect 9739 2692 9763 2694
rect 9819 2692 9825 2694
rect 9517 2683 9825 2692
rect 10796 2446 10824 4422
rect 11230 4380 11538 4389
rect 11230 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11396 4380
rect 11452 4378 11476 4380
rect 11532 4378 11538 4380
rect 11292 4326 11294 4378
rect 11474 4326 11476 4378
rect 11230 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11396 4326
rect 11452 4324 11476 4326
rect 11532 4324 11538 4326
rect 11230 4315 11538 4324
rect 14657 4380 14965 4389
rect 14657 4378 14663 4380
rect 14719 4378 14743 4380
rect 14799 4378 14823 4380
rect 14879 4378 14903 4380
rect 14959 4378 14965 4380
rect 14719 4326 14721 4378
rect 14901 4326 14903 4378
rect 14657 4324 14663 4326
rect 14719 4324 14743 4326
rect 14799 4324 14823 4326
rect 14879 4324 14903 4326
rect 14959 4324 14965 4326
rect 14657 4315 14965 4324
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 12944 3836 13252 3845
rect 12944 3834 12950 3836
rect 13006 3834 13030 3836
rect 13086 3834 13110 3836
rect 13166 3834 13190 3836
rect 13246 3834 13252 3836
rect 13006 3782 13008 3834
rect 13188 3782 13190 3834
rect 12944 3780 12950 3782
rect 13006 3780 13030 3782
rect 13086 3780 13110 3782
rect 13166 3780 13190 3782
rect 13246 3780 13252 3782
rect 12944 3771 13252 3780
rect 11230 3292 11538 3301
rect 11230 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11396 3292
rect 11452 3290 11476 3292
rect 11532 3290 11538 3292
rect 11292 3238 11294 3290
rect 11474 3238 11476 3290
rect 11230 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11396 3238
rect 11452 3236 11476 3238
rect 11532 3236 11538 3238
rect 11230 3227 11538 3236
rect 12944 2748 13252 2757
rect 12944 2746 12950 2748
rect 13006 2746 13030 2748
rect 13086 2746 13110 2748
rect 13166 2746 13190 2748
rect 13246 2746 13252 2748
rect 13006 2694 13008 2746
rect 13188 2694 13190 2746
rect 12944 2692 12950 2694
rect 13006 2692 13030 2694
rect 13086 2692 13110 2694
rect 13166 2692 13190 2694
rect 13246 2692 13252 2694
rect 12944 2683 13252 2692
rect 13464 2446 13492 4218
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 14016 3058 14044 3334
rect 14657 3292 14965 3301
rect 14657 3290 14663 3292
rect 14719 3290 14743 3292
rect 14799 3290 14823 3292
rect 14879 3290 14903 3292
rect 14959 3290 14965 3292
rect 14719 3238 14721 3290
rect 14901 3238 14903 3290
rect 14657 3236 14663 3238
rect 14719 3236 14743 3238
rect 14799 3236 14823 3238
rect 14879 3236 14903 3238
rect 14959 3236 14965 3238
rect 14657 3227 14965 3236
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 1032 2304 1084 2310
rect 1032 2246 1084 2252
rect 2412 2304 2464 2310
rect 2412 2246 2464 2252
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 1044 800 1072 2246
rect 2424 800 2452 2246
rect 3804 800 3832 2246
rect 4376 2204 4684 2213
rect 4376 2202 4382 2204
rect 4438 2202 4462 2204
rect 4518 2202 4542 2204
rect 4598 2202 4622 2204
rect 4678 2202 4684 2204
rect 4438 2150 4440 2202
rect 4620 2150 4622 2202
rect 4376 2148 4382 2150
rect 4438 2148 4462 2150
rect 4518 2148 4542 2150
rect 4598 2148 4622 2150
rect 4678 2148 4684 2150
rect 4376 2139 4684 2148
rect 5184 800 5212 2246
rect 6564 800 6592 2246
rect 7803 2204 8111 2213
rect 7803 2202 7809 2204
rect 7865 2202 7889 2204
rect 7945 2202 7969 2204
rect 8025 2202 8049 2204
rect 8105 2202 8111 2204
rect 7865 2150 7867 2202
rect 8047 2150 8049 2202
rect 7803 2148 7809 2150
rect 7865 2148 7889 2150
rect 7945 2148 7969 2150
rect 8025 2148 8049 2150
rect 8105 2148 8111 2150
rect 7803 2139 8111 2148
rect 7944 870 8064 898
rect 7944 800 7972 870
rect 1030 0 1086 800
rect 2410 0 2466 800
rect 3790 0 3846 800
rect 5170 0 5226 800
rect 6550 0 6606 800
rect 7930 0 7986 800
rect 8036 762 8064 870
rect 8220 762 8248 2246
rect 9324 800 9352 2246
rect 10704 800 10732 2246
rect 11230 2204 11538 2213
rect 11230 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11396 2204
rect 11452 2202 11476 2204
rect 11532 2202 11538 2204
rect 11292 2150 11294 2202
rect 11474 2150 11476 2202
rect 11230 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11396 2150
rect 11452 2148 11476 2150
rect 11532 2148 11538 2150
rect 11230 2139 11538 2148
rect 12084 800 12112 2246
rect 13464 800 13492 2246
rect 8036 734 8248 762
rect 9310 0 9366 800
rect 10690 0 10746 800
rect 12070 0 12126 800
rect 13450 0 13506 800
rect 14568 762 14596 2790
rect 14657 2204 14965 2213
rect 14657 2202 14663 2204
rect 14719 2202 14743 2204
rect 14799 2202 14823 2204
rect 14879 2202 14903 2204
rect 14959 2202 14965 2204
rect 14719 2150 14721 2202
rect 14901 2150 14903 2202
rect 14657 2148 14663 2150
rect 14719 2148 14743 2150
rect 14799 2148 14823 2150
rect 14879 2148 14903 2150
rect 14959 2148 14965 2150
rect 14657 2139 14965 2148
rect 14752 870 14872 898
rect 14752 762 14780 870
rect 14844 800 14872 870
rect 14568 734 14780 762
rect 14830 0 14886 800
<< via2 >>
rect 2669 6010 2725 6012
rect 2749 6010 2805 6012
rect 2829 6010 2885 6012
rect 2909 6010 2965 6012
rect 2669 5958 2715 6010
rect 2715 5958 2725 6010
rect 2749 5958 2779 6010
rect 2779 5958 2791 6010
rect 2791 5958 2805 6010
rect 2829 5958 2843 6010
rect 2843 5958 2855 6010
rect 2855 5958 2885 6010
rect 2909 5958 2919 6010
rect 2919 5958 2965 6010
rect 2669 5956 2725 5958
rect 2749 5956 2805 5958
rect 2829 5956 2885 5958
rect 2909 5956 2965 5958
rect 4382 6554 4438 6556
rect 4462 6554 4518 6556
rect 4542 6554 4598 6556
rect 4622 6554 4678 6556
rect 4382 6502 4428 6554
rect 4428 6502 4438 6554
rect 4462 6502 4492 6554
rect 4492 6502 4504 6554
rect 4504 6502 4518 6554
rect 4542 6502 4556 6554
rect 4556 6502 4568 6554
rect 4568 6502 4598 6554
rect 4622 6502 4632 6554
rect 4632 6502 4678 6554
rect 4382 6500 4438 6502
rect 4462 6500 4518 6502
rect 4542 6500 4598 6502
rect 4622 6500 4678 6502
rect 7809 6554 7865 6556
rect 7889 6554 7945 6556
rect 7969 6554 8025 6556
rect 8049 6554 8105 6556
rect 7809 6502 7855 6554
rect 7855 6502 7865 6554
rect 7889 6502 7919 6554
rect 7919 6502 7931 6554
rect 7931 6502 7945 6554
rect 7969 6502 7983 6554
rect 7983 6502 7995 6554
rect 7995 6502 8025 6554
rect 8049 6502 8059 6554
rect 8059 6502 8105 6554
rect 7809 6500 7865 6502
rect 7889 6500 7945 6502
rect 7969 6500 8025 6502
rect 8049 6500 8105 6502
rect 2669 4922 2725 4924
rect 2749 4922 2805 4924
rect 2829 4922 2885 4924
rect 2909 4922 2965 4924
rect 2669 4870 2715 4922
rect 2715 4870 2725 4922
rect 2749 4870 2779 4922
rect 2779 4870 2791 4922
rect 2791 4870 2805 4922
rect 2829 4870 2843 4922
rect 2843 4870 2855 4922
rect 2855 4870 2885 4922
rect 2909 4870 2919 4922
rect 2919 4870 2965 4922
rect 2669 4868 2725 4870
rect 2749 4868 2805 4870
rect 2829 4868 2885 4870
rect 2909 4868 2965 4870
rect 4382 5466 4438 5468
rect 4462 5466 4518 5468
rect 4542 5466 4598 5468
rect 4622 5466 4678 5468
rect 4382 5414 4428 5466
rect 4428 5414 4438 5466
rect 4462 5414 4492 5466
rect 4492 5414 4504 5466
rect 4504 5414 4518 5466
rect 4542 5414 4556 5466
rect 4556 5414 4568 5466
rect 4568 5414 4598 5466
rect 4622 5414 4632 5466
rect 4632 5414 4678 5466
rect 4382 5412 4438 5414
rect 4462 5412 4518 5414
rect 4542 5412 4598 5414
rect 4622 5412 4678 5414
rect 4382 4378 4438 4380
rect 4462 4378 4518 4380
rect 4542 4378 4598 4380
rect 4622 4378 4678 4380
rect 4382 4326 4428 4378
rect 4428 4326 4438 4378
rect 4462 4326 4492 4378
rect 4492 4326 4504 4378
rect 4504 4326 4518 4378
rect 4542 4326 4556 4378
rect 4556 4326 4568 4378
rect 4568 4326 4598 4378
rect 4622 4326 4632 4378
rect 4632 4326 4678 4378
rect 4382 4324 4438 4326
rect 4462 4324 4518 4326
rect 4542 4324 4598 4326
rect 4622 4324 4678 4326
rect 2669 3834 2725 3836
rect 2749 3834 2805 3836
rect 2829 3834 2885 3836
rect 2909 3834 2965 3836
rect 2669 3782 2715 3834
rect 2715 3782 2725 3834
rect 2749 3782 2779 3834
rect 2779 3782 2791 3834
rect 2791 3782 2805 3834
rect 2829 3782 2843 3834
rect 2843 3782 2855 3834
rect 2855 3782 2885 3834
rect 2909 3782 2919 3834
rect 2919 3782 2965 3834
rect 2669 3780 2725 3782
rect 2749 3780 2805 3782
rect 2829 3780 2885 3782
rect 2909 3780 2965 3782
rect 2669 2746 2725 2748
rect 2749 2746 2805 2748
rect 2829 2746 2885 2748
rect 2909 2746 2965 2748
rect 2669 2694 2715 2746
rect 2715 2694 2725 2746
rect 2749 2694 2779 2746
rect 2779 2694 2791 2746
rect 2791 2694 2805 2746
rect 2829 2694 2843 2746
rect 2843 2694 2855 2746
rect 2855 2694 2885 2746
rect 2909 2694 2919 2746
rect 2919 2694 2965 2746
rect 2669 2692 2725 2694
rect 2749 2692 2805 2694
rect 2829 2692 2885 2694
rect 2909 2692 2965 2694
rect 4382 3290 4438 3292
rect 4462 3290 4518 3292
rect 4542 3290 4598 3292
rect 4622 3290 4678 3292
rect 4382 3238 4428 3290
rect 4428 3238 4438 3290
rect 4462 3238 4492 3290
rect 4492 3238 4504 3290
rect 4504 3238 4518 3290
rect 4542 3238 4556 3290
rect 4556 3238 4568 3290
rect 4568 3238 4598 3290
rect 4622 3238 4632 3290
rect 4632 3238 4678 3290
rect 4382 3236 4438 3238
rect 4462 3236 4518 3238
rect 4542 3236 4598 3238
rect 4622 3236 4678 3238
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6096 5958 6142 6010
rect 6142 5958 6152 6010
rect 6176 5958 6206 6010
rect 6206 5958 6218 6010
rect 6218 5958 6232 6010
rect 6256 5958 6270 6010
rect 6270 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6096 4870 6142 4922
rect 6142 4870 6152 4922
rect 6176 4870 6206 4922
rect 6206 4870 6218 4922
rect 6218 4870 6232 4922
rect 6256 4870 6270 4922
rect 6270 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11396 6554 11452 6556
rect 11476 6554 11532 6556
rect 11236 6502 11282 6554
rect 11282 6502 11292 6554
rect 11316 6502 11346 6554
rect 11346 6502 11358 6554
rect 11358 6502 11372 6554
rect 11396 6502 11410 6554
rect 11410 6502 11422 6554
rect 11422 6502 11452 6554
rect 11476 6502 11486 6554
rect 11486 6502 11532 6554
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11396 6500 11452 6502
rect 11476 6500 11532 6502
rect 14663 6554 14719 6556
rect 14743 6554 14799 6556
rect 14823 6554 14879 6556
rect 14903 6554 14959 6556
rect 14663 6502 14709 6554
rect 14709 6502 14719 6554
rect 14743 6502 14773 6554
rect 14773 6502 14785 6554
rect 14785 6502 14799 6554
rect 14823 6502 14837 6554
rect 14837 6502 14849 6554
rect 14849 6502 14879 6554
rect 14903 6502 14913 6554
rect 14913 6502 14959 6554
rect 14663 6500 14719 6502
rect 14743 6500 14799 6502
rect 14823 6500 14879 6502
rect 14903 6500 14959 6502
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6096 3782 6142 3834
rect 6142 3782 6152 3834
rect 6176 3782 6206 3834
rect 6206 3782 6218 3834
rect 6218 3782 6232 3834
rect 6256 3782 6270 3834
rect 6270 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6096 2694 6142 2746
rect 6142 2694 6152 2746
rect 6176 2694 6206 2746
rect 6206 2694 6218 2746
rect 6218 2694 6232 2746
rect 6256 2694 6270 2746
rect 6270 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 9523 6010 9579 6012
rect 9603 6010 9659 6012
rect 9683 6010 9739 6012
rect 9763 6010 9819 6012
rect 9523 5958 9569 6010
rect 9569 5958 9579 6010
rect 9603 5958 9633 6010
rect 9633 5958 9645 6010
rect 9645 5958 9659 6010
rect 9683 5958 9697 6010
rect 9697 5958 9709 6010
rect 9709 5958 9739 6010
rect 9763 5958 9773 6010
rect 9773 5958 9819 6010
rect 9523 5956 9579 5958
rect 9603 5956 9659 5958
rect 9683 5956 9739 5958
rect 9763 5956 9819 5958
rect 12950 6010 13006 6012
rect 13030 6010 13086 6012
rect 13110 6010 13166 6012
rect 13190 6010 13246 6012
rect 12950 5958 12996 6010
rect 12996 5958 13006 6010
rect 13030 5958 13060 6010
rect 13060 5958 13072 6010
rect 13072 5958 13086 6010
rect 13110 5958 13124 6010
rect 13124 5958 13136 6010
rect 13136 5958 13166 6010
rect 13190 5958 13200 6010
rect 13200 5958 13246 6010
rect 12950 5956 13006 5958
rect 13030 5956 13086 5958
rect 13110 5956 13166 5958
rect 13190 5956 13246 5958
rect 7809 5466 7865 5468
rect 7889 5466 7945 5468
rect 7969 5466 8025 5468
rect 8049 5466 8105 5468
rect 7809 5414 7855 5466
rect 7855 5414 7865 5466
rect 7889 5414 7919 5466
rect 7919 5414 7931 5466
rect 7931 5414 7945 5466
rect 7969 5414 7983 5466
rect 7983 5414 7995 5466
rect 7995 5414 8025 5466
rect 8049 5414 8059 5466
rect 8059 5414 8105 5466
rect 7809 5412 7865 5414
rect 7889 5412 7945 5414
rect 7969 5412 8025 5414
rect 8049 5412 8105 5414
rect 7809 4378 7865 4380
rect 7889 4378 7945 4380
rect 7969 4378 8025 4380
rect 8049 4378 8105 4380
rect 7809 4326 7855 4378
rect 7855 4326 7865 4378
rect 7889 4326 7919 4378
rect 7919 4326 7931 4378
rect 7931 4326 7945 4378
rect 7969 4326 7983 4378
rect 7983 4326 7995 4378
rect 7995 4326 8025 4378
rect 8049 4326 8059 4378
rect 8059 4326 8105 4378
rect 7809 4324 7865 4326
rect 7889 4324 7945 4326
rect 7969 4324 8025 4326
rect 8049 4324 8105 4326
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11396 5466 11452 5468
rect 11476 5466 11532 5468
rect 11236 5414 11282 5466
rect 11282 5414 11292 5466
rect 11316 5414 11346 5466
rect 11346 5414 11358 5466
rect 11358 5414 11372 5466
rect 11396 5414 11410 5466
rect 11410 5414 11422 5466
rect 11422 5414 11452 5466
rect 11476 5414 11486 5466
rect 11486 5414 11532 5466
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11396 5412 11452 5414
rect 11476 5412 11532 5414
rect 14663 5466 14719 5468
rect 14743 5466 14799 5468
rect 14823 5466 14879 5468
rect 14903 5466 14959 5468
rect 14663 5414 14709 5466
rect 14709 5414 14719 5466
rect 14743 5414 14773 5466
rect 14773 5414 14785 5466
rect 14785 5414 14799 5466
rect 14823 5414 14837 5466
rect 14837 5414 14849 5466
rect 14849 5414 14879 5466
rect 14903 5414 14913 5466
rect 14913 5414 14959 5466
rect 14663 5412 14719 5414
rect 14743 5412 14799 5414
rect 14823 5412 14879 5414
rect 14903 5412 14959 5414
rect 9523 4922 9579 4924
rect 9603 4922 9659 4924
rect 9683 4922 9739 4924
rect 9763 4922 9819 4924
rect 9523 4870 9569 4922
rect 9569 4870 9579 4922
rect 9603 4870 9633 4922
rect 9633 4870 9645 4922
rect 9645 4870 9659 4922
rect 9683 4870 9697 4922
rect 9697 4870 9709 4922
rect 9709 4870 9739 4922
rect 9763 4870 9773 4922
rect 9773 4870 9819 4922
rect 9523 4868 9579 4870
rect 9603 4868 9659 4870
rect 9683 4868 9739 4870
rect 9763 4868 9819 4870
rect 12950 4922 13006 4924
rect 13030 4922 13086 4924
rect 13110 4922 13166 4924
rect 13190 4922 13246 4924
rect 12950 4870 12996 4922
rect 12996 4870 13006 4922
rect 13030 4870 13060 4922
rect 13060 4870 13072 4922
rect 13072 4870 13086 4922
rect 13110 4870 13124 4922
rect 13124 4870 13136 4922
rect 13136 4870 13166 4922
rect 13190 4870 13200 4922
rect 13200 4870 13246 4922
rect 12950 4868 13006 4870
rect 13030 4868 13086 4870
rect 13110 4868 13166 4870
rect 13190 4868 13246 4870
rect 7809 3290 7865 3292
rect 7889 3290 7945 3292
rect 7969 3290 8025 3292
rect 8049 3290 8105 3292
rect 7809 3238 7855 3290
rect 7855 3238 7865 3290
rect 7889 3238 7919 3290
rect 7919 3238 7931 3290
rect 7931 3238 7945 3290
rect 7969 3238 7983 3290
rect 7983 3238 7995 3290
rect 7995 3238 8025 3290
rect 8049 3238 8059 3290
rect 8059 3238 8105 3290
rect 7809 3236 7865 3238
rect 7889 3236 7945 3238
rect 7969 3236 8025 3238
rect 8049 3236 8105 3238
rect 9523 3834 9579 3836
rect 9603 3834 9659 3836
rect 9683 3834 9739 3836
rect 9763 3834 9819 3836
rect 9523 3782 9569 3834
rect 9569 3782 9579 3834
rect 9603 3782 9633 3834
rect 9633 3782 9645 3834
rect 9645 3782 9659 3834
rect 9683 3782 9697 3834
rect 9697 3782 9709 3834
rect 9709 3782 9739 3834
rect 9763 3782 9773 3834
rect 9773 3782 9819 3834
rect 9523 3780 9579 3782
rect 9603 3780 9659 3782
rect 9683 3780 9739 3782
rect 9763 3780 9819 3782
rect 9523 2746 9579 2748
rect 9603 2746 9659 2748
rect 9683 2746 9739 2748
rect 9763 2746 9819 2748
rect 9523 2694 9569 2746
rect 9569 2694 9579 2746
rect 9603 2694 9633 2746
rect 9633 2694 9645 2746
rect 9645 2694 9659 2746
rect 9683 2694 9697 2746
rect 9697 2694 9709 2746
rect 9709 2694 9739 2746
rect 9763 2694 9773 2746
rect 9773 2694 9819 2746
rect 9523 2692 9579 2694
rect 9603 2692 9659 2694
rect 9683 2692 9739 2694
rect 9763 2692 9819 2694
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11396 4378 11452 4380
rect 11476 4378 11532 4380
rect 11236 4326 11282 4378
rect 11282 4326 11292 4378
rect 11316 4326 11346 4378
rect 11346 4326 11358 4378
rect 11358 4326 11372 4378
rect 11396 4326 11410 4378
rect 11410 4326 11422 4378
rect 11422 4326 11452 4378
rect 11476 4326 11486 4378
rect 11486 4326 11532 4378
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 11396 4324 11452 4326
rect 11476 4324 11532 4326
rect 14663 4378 14719 4380
rect 14743 4378 14799 4380
rect 14823 4378 14879 4380
rect 14903 4378 14959 4380
rect 14663 4326 14709 4378
rect 14709 4326 14719 4378
rect 14743 4326 14773 4378
rect 14773 4326 14785 4378
rect 14785 4326 14799 4378
rect 14823 4326 14837 4378
rect 14837 4326 14849 4378
rect 14849 4326 14879 4378
rect 14903 4326 14913 4378
rect 14913 4326 14959 4378
rect 14663 4324 14719 4326
rect 14743 4324 14799 4326
rect 14823 4324 14879 4326
rect 14903 4324 14959 4326
rect 12950 3834 13006 3836
rect 13030 3834 13086 3836
rect 13110 3834 13166 3836
rect 13190 3834 13246 3836
rect 12950 3782 12996 3834
rect 12996 3782 13006 3834
rect 13030 3782 13060 3834
rect 13060 3782 13072 3834
rect 13072 3782 13086 3834
rect 13110 3782 13124 3834
rect 13124 3782 13136 3834
rect 13136 3782 13166 3834
rect 13190 3782 13200 3834
rect 13200 3782 13246 3834
rect 12950 3780 13006 3782
rect 13030 3780 13086 3782
rect 13110 3780 13166 3782
rect 13190 3780 13246 3782
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11396 3290 11452 3292
rect 11476 3290 11532 3292
rect 11236 3238 11282 3290
rect 11282 3238 11292 3290
rect 11316 3238 11346 3290
rect 11346 3238 11358 3290
rect 11358 3238 11372 3290
rect 11396 3238 11410 3290
rect 11410 3238 11422 3290
rect 11422 3238 11452 3290
rect 11476 3238 11486 3290
rect 11486 3238 11532 3290
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11396 3236 11452 3238
rect 11476 3236 11532 3238
rect 12950 2746 13006 2748
rect 13030 2746 13086 2748
rect 13110 2746 13166 2748
rect 13190 2746 13246 2748
rect 12950 2694 12996 2746
rect 12996 2694 13006 2746
rect 13030 2694 13060 2746
rect 13060 2694 13072 2746
rect 13072 2694 13086 2746
rect 13110 2694 13124 2746
rect 13124 2694 13136 2746
rect 13136 2694 13166 2746
rect 13190 2694 13200 2746
rect 13200 2694 13246 2746
rect 12950 2692 13006 2694
rect 13030 2692 13086 2694
rect 13110 2692 13166 2694
rect 13190 2692 13246 2694
rect 14663 3290 14719 3292
rect 14743 3290 14799 3292
rect 14823 3290 14879 3292
rect 14903 3290 14959 3292
rect 14663 3238 14709 3290
rect 14709 3238 14719 3290
rect 14743 3238 14773 3290
rect 14773 3238 14785 3290
rect 14785 3238 14799 3290
rect 14823 3238 14837 3290
rect 14837 3238 14849 3290
rect 14849 3238 14879 3290
rect 14903 3238 14913 3290
rect 14913 3238 14959 3290
rect 14663 3236 14719 3238
rect 14743 3236 14799 3238
rect 14823 3236 14879 3238
rect 14903 3236 14959 3238
rect 4382 2202 4438 2204
rect 4462 2202 4518 2204
rect 4542 2202 4598 2204
rect 4622 2202 4678 2204
rect 4382 2150 4428 2202
rect 4428 2150 4438 2202
rect 4462 2150 4492 2202
rect 4492 2150 4504 2202
rect 4504 2150 4518 2202
rect 4542 2150 4556 2202
rect 4556 2150 4568 2202
rect 4568 2150 4598 2202
rect 4622 2150 4632 2202
rect 4632 2150 4678 2202
rect 4382 2148 4438 2150
rect 4462 2148 4518 2150
rect 4542 2148 4598 2150
rect 4622 2148 4678 2150
rect 7809 2202 7865 2204
rect 7889 2202 7945 2204
rect 7969 2202 8025 2204
rect 8049 2202 8105 2204
rect 7809 2150 7855 2202
rect 7855 2150 7865 2202
rect 7889 2150 7919 2202
rect 7919 2150 7931 2202
rect 7931 2150 7945 2202
rect 7969 2150 7983 2202
rect 7983 2150 7995 2202
rect 7995 2150 8025 2202
rect 8049 2150 8059 2202
rect 8059 2150 8105 2202
rect 7809 2148 7865 2150
rect 7889 2148 7945 2150
rect 7969 2148 8025 2150
rect 8049 2148 8105 2150
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11396 2202 11452 2204
rect 11476 2202 11532 2204
rect 11236 2150 11282 2202
rect 11282 2150 11292 2202
rect 11316 2150 11346 2202
rect 11346 2150 11358 2202
rect 11358 2150 11372 2202
rect 11396 2150 11410 2202
rect 11410 2150 11422 2202
rect 11422 2150 11452 2202
rect 11476 2150 11486 2202
rect 11486 2150 11532 2202
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 11396 2148 11452 2150
rect 11476 2148 11532 2150
rect 14663 2202 14719 2204
rect 14743 2202 14799 2204
rect 14823 2202 14879 2204
rect 14903 2202 14959 2204
rect 14663 2150 14709 2202
rect 14709 2150 14719 2202
rect 14743 2150 14773 2202
rect 14773 2150 14785 2202
rect 14785 2150 14799 2202
rect 14823 2150 14837 2202
rect 14837 2150 14849 2202
rect 14849 2150 14879 2202
rect 14903 2150 14913 2202
rect 14913 2150 14959 2202
rect 14663 2148 14719 2150
rect 14743 2148 14799 2150
rect 14823 2148 14879 2150
rect 14903 2148 14959 2150
<< metal3 >>
rect 4372 6560 4688 6561
rect 4372 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4688 6560
rect 4372 6495 4688 6496
rect 7799 6560 8115 6561
rect 7799 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8115 6560
rect 7799 6495 8115 6496
rect 11226 6560 11542 6561
rect 11226 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11542 6560
rect 11226 6495 11542 6496
rect 14653 6560 14969 6561
rect 14653 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14969 6560
rect 14653 6495 14969 6496
rect 2659 6016 2975 6017
rect 2659 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2975 6016
rect 2659 5951 2975 5952
rect 6086 6016 6402 6017
rect 6086 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6402 6016
rect 6086 5951 6402 5952
rect 9513 6016 9829 6017
rect 9513 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9829 6016
rect 9513 5951 9829 5952
rect 12940 6016 13256 6017
rect 12940 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13256 6016
rect 12940 5951 13256 5952
rect 4372 5472 4688 5473
rect 4372 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4688 5472
rect 4372 5407 4688 5408
rect 7799 5472 8115 5473
rect 7799 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8115 5472
rect 7799 5407 8115 5408
rect 11226 5472 11542 5473
rect 11226 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11542 5472
rect 11226 5407 11542 5408
rect 14653 5472 14969 5473
rect 14653 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14969 5472
rect 14653 5407 14969 5408
rect 2659 4928 2975 4929
rect 2659 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2975 4928
rect 2659 4863 2975 4864
rect 6086 4928 6402 4929
rect 6086 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6402 4928
rect 6086 4863 6402 4864
rect 9513 4928 9829 4929
rect 9513 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9829 4928
rect 9513 4863 9829 4864
rect 12940 4928 13256 4929
rect 12940 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13256 4928
rect 12940 4863 13256 4864
rect 4372 4384 4688 4385
rect 4372 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4688 4384
rect 4372 4319 4688 4320
rect 7799 4384 8115 4385
rect 7799 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8115 4384
rect 7799 4319 8115 4320
rect 11226 4384 11542 4385
rect 11226 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11542 4384
rect 11226 4319 11542 4320
rect 14653 4384 14969 4385
rect 14653 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14969 4384
rect 14653 4319 14969 4320
rect 2659 3840 2975 3841
rect 2659 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2975 3840
rect 2659 3775 2975 3776
rect 6086 3840 6402 3841
rect 6086 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6402 3840
rect 6086 3775 6402 3776
rect 9513 3840 9829 3841
rect 9513 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9829 3840
rect 9513 3775 9829 3776
rect 12940 3840 13256 3841
rect 12940 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13256 3840
rect 12940 3775 13256 3776
rect 4372 3296 4688 3297
rect 4372 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4688 3296
rect 4372 3231 4688 3232
rect 7799 3296 8115 3297
rect 7799 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8115 3296
rect 7799 3231 8115 3232
rect 11226 3296 11542 3297
rect 11226 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11542 3296
rect 11226 3231 11542 3232
rect 14653 3296 14969 3297
rect 14653 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14969 3296
rect 14653 3231 14969 3232
rect 2659 2752 2975 2753
rect 2659 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2975 2752
rect 2659 2687 2975 2688
rect 6086 2752 6402 2753
rect 6086 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6402 2752
rect 6086 2687 6402 2688
rect 9513 2752 9829 2753
rect 9513 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9829 2752
rect 9513 2687 9829 2688
rect 12940 2752 13256 2753
rect 12940 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13256 2752
rect 12940 2687 13256 2688
rect 4372 2208 4688 2209
rect 4372 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4688 2208
rect 4372 2143 4688 2144
rect 7799 2208 8115 2209
rect 7799 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8115 2208
rect 7799 2143 8115 2144
rect 11226 2208 11542 2209
rect 11226 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11542 2208
rect 11226 2143 11542 2144
rect 14653 2208 14969 2209
rect 14653 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14969 2208
rect 14653 2143 14969 2144
<< via3 >>
rect 4378 6556 4442 6560
rect 4378 6500 4382 6556
rect 4382 6500 4438 6556
rect 4438 6500 4442 6556
rect 4378 6496 4442 6500
rect 4458 6556 4522 6560
rect 4458 6500 4462 6556
rect 4462 6500 4518 6556
rect 4518 6500 4522 6556
rect 4458 6496 4522 6500
rect 4538 6556 4602 6560
rect 4538 6500 4542 6556
rect 4542 6500 4598 6556
rect 4598 6500 4602 6556
rect 4538 6496 4602 6500
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 7805 6556 7869 6560
rect 7805 6500 7809 6556
rect 7809 6500 7865 6556
rect 7865 6500 7869 6556
rect 7805 6496 7869 6500
rect 7885 6556 7949 6560
rect 7885 6500 7889 6556
rect 7889 6500 7945 6556
rect 7945 6500 7949 6556
rect 7885 6496 7949 6500
rect 7965 6556 8029 6560
rect 7965 6500 7969 6556
rect 7969 6500 8025 6556
rect 8025 6500 8029 6556
rect 7965 6496 8029 6500
rect 8045 6556 8109 6560
rect 8045 6500 8049 6556
rect 8049 6500 8105 6556
rect 8105 6500 8109 6556
rect 8045 6496 8109 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 11392 6556 11456 6560
rect 11392 6500 11396 6556
rect 11396 6500 11452 6556
rect 11452 6500 11456 6556
rect 11392 6496 11456 6500
rect 11472 6556 11536 6560
rect 11472 6500 11476 6556
rect 11476 6500 11532 6556
rect 11532 6500 11536 6556
rect 11472 6496 11536 6500
rect 14659 6556 14723 6560
rect 14659 6500 14663 6556
rect 14663 6500 14719 6556
rect 14719 6500 14723 6556
rect 14659 6496 14723 6500
rect 14739 6556 14803 6560
rect 14739 6500 14743 6556
rect 14743 6500 14799 6556
rect 14799 6500 14803 6556
rect 14739 6496 14803 6500
rect 14819 6556 14883 6560
rect 14819 6500 14823 6556
rect 14823 6500 14879 6556
rect 14879 6500 14883 6556
rect 14819 6496 14883 6500
rect 14899 6556 14963 6560
rect 14899 6500 14903 6556
rect 14903 6500 14959 6556
rect 14959 6500 14963 6556
rect 14899 6496 14963 6500
rect 2665 6012 2729 6016
rect 2665 5956 2669 6012
rect 2669 5956 2725 6012
rect 2725 5956 2729 6012
rect 2665 5952 2729 5956
rect 2745 6012 2809 6016
rect 2745 5956 2749 6012
rect 2749 5956 2805 6012
rect 2805 5956 2809 6012
rect 2745 5952 2809 5956
rect 2825 6012 2889 6016
rect 2825 5956 2829 6012
rect 2829 5956 2885 6012
rect 2885 5956 2889 6012
rect 2825 5952 2889 5956
rect 2905 6012 2969 6016
rect 2905 5956 2909 6012
rect 2909 5956 2965 6012
rect 2965 5956 2969 6012
rect 2905 5952 2969 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 9519 6012 9583 6016
rect 9519 5956 9523 6012
rect 9523 5956 9579 6012
rect 9579 5956 9583 6012
rect 9519 5952 9583 5956
rect 9599 6012 9663 6016
rect 9599 5956 9603 6012
rect 9603 5956 9659 6012
rect 9659 5956 9663 6012
rect 9599 5952 9663 5956
rect 9679 6012 9743 6016
rect 9679 5956 9683 6012
rect 9683 5956 9739 6012
rect 9739 5956 9743 6012
rect 9679 5952 9743 5956
rect 9759 6012 9823 6016
rect 9759 5956 9763 6012
rect 9763 5956 9819 6012
rect 9819 5956 9823 6012
rect 9759 5952 9823 5956
rect 12946 6012 13010 6016
rect 12946 5956 12950 6012
rect 12950 5956 13006 6012
rect 13006 5956 13010 6012
rect 12946 5952 13010 5956
rect 13026 6012 13090 6016
rect 13026 5956 13030 6012
rect 13030 5956 13086 6012
rect 13086 5956 13090 6012
rect 13026 5952 13090 5956
rect 13106 6012 13170 6016
rect 13106 5956 13110 6012
rect 13110 5956 13166 6012
rect 13166 5956 13170 6012
rect 13106 5952 13170 5956
rect 13186 6012 13250 6016
rect 13186 5956 13190 6012
rect 13190 5956 13246 6012
rect 13246 5956 13250 6012
rect 13186 5952 13250 5956
rect 4378 5468 4442 5472
rect 4378 5412 4382 5468
rect 4382 5412 4438 5468
rect 4438 5412 4442 5468
rect 4378 5408 4442 5412
rect 4458 5468 4522 5472
rect 4458 5412 4462 5468
rect 4462 5412 4518 5468
rect 4518 5412 4522 5468
rect 4458 5408 4522 5412
rect 4538 5468 4602 5472
rect 4538 5412 4542 5468
rect 4542 5412 4598 5468
rect 4598 5412 4602 5468
rect 4538 5408 4602 5412
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 7805 5468 7869 5472
rect 7805 5412 7809 5468
rect 7809 5412 7865 5468
rect 7865 5412 7869 5468
rect 7805 5408 7869 5412
rect 7885 5468 7949 5472
rect 7885 5412 7889 5468
rect 7889 5412 7945 5468
rect 7945 5412 7949 5468
rect 7885 5408 7949 5412
rect 7965 5468 8029 5472
rect 7965 5412 7969 5468
rect 7969 5412 8025 5468
rect 8025 5412 8029 5468
rect 7965 5408 8029 5412
rect 8045 5468 8109 5472
rect 8045 5412 8049 5468
rect 8049 5412 8105 5468
rect 8105 5412 8109 5468
rect 8045 5408 8109 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 11392 5468 11456 5472
rect 11392 5412 11396 5468
rect 11396 5412 11452 5468
rect 11452 5412 11456 5468
rect 11392 5408 11456 5412
rect 11472 5468 11536 5472
rect 11472 5412 11476 5468
rect 11476 5412 11532 5468
rect 11532 5412 11536 5468
rect 11472 5408 11536 5412
rect 14659 5468 14723 5472
rect 14659 5412 14663 5468
rect 14663 5412 14719 5468
rect 14719 5412 14723 5468
rect 14659 5408 14723 5412
rect 14739 5468 14803 5472
rect 14739 5412 14743 5468
rect 14743 5412 14799 5468
rect 14799 5412 14803 5468
rect 14739 5408 14803 5412
rect 14819 5468 14883 5472
rect 14819 5412 14823 5468
rect 14823 5412 14879 5468
rect 14879 5412 14883 5468
rect 14819 5408 14883 5412
rect 14899 5468 14963 5472
rect 14899 5412 14903 5468
rect 14903 5412 14959 5468
rect 14959 5412 14963 5468
rect 14899 5408 14963 5412
rect 2665 4924 2729 4928
rect 2665 4868 2669 4924
rect 2669 4868 2725 4924
rect 2725 4868 2729 4924
rect 2665 4864 2729 4868
rect 2745 4924 2809 4928
rect 2745 4868 2749 4924
rect 2749 4868 2805 4924
rect 2805 4868 2809 4924
rect 2745 4864 2809 4868
rect 2825 4924 2889 4928
rect 2825 4868 2829 4924
rect 2829 4868 2885 4924
rect 2885 4868 2889 4924
rect 2825 4864 2889 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 9519 4924 9583 4928
rect 9519 4868 9523 4924
rect 9523 4868 9579 4924
rect 9579 4868 9583 4924
rect 9519 4864 9583 4868
rect 9599 4924 9663 4928
rect 9599 4868 9603 4924
rect 9603 4868 9659 4924
rect 9659 4868 9663 4924
rect 9599 4864 9663 4868
rect 9679 4924 9743 4928
rect 9679 4868 9683 4924
rect 9683 4868 9739 4924
rect 9739 4868 9743 4924
rect 9679 4864 9743 4868
rect 9759 4924 9823 4928
rect 9759 4868 9763 4924
rect 9763 4868 9819 4924
rect 9819 4868 9823 4924
rect 9759 4864 9823 4868
rect 12946 4924 13010 4928
rect 12946 4868 12950 4924
rect 12950 4868 13006 4924
rect 13006 4868 13010 4924
rect 12946 4864 13010 4868
rect 13026 4924 13090 4928
rect 13026 4868 13030 4924
rect 13030 4868 13086 4924
rect 13086 4868 13090 4924
rect 13026 4864 13090 4868
rect 13106 4924 13170 4928
rect 13106 4868 13110 4924
rect 13110 4868 13166 4924
rect 13166 4868 13170 4924
rect 13106 4864 13170 4868
rect 13186 4924 13250 4928
rect 13186 4868 13190 4924
rect 13190 4868 13246 4924
rect 13246 4868 13250 4924
rect 13186 4864 13250 4868
rect 4378 4380 4442 4384
rect 4378 4324 4382 4380
rect 4382 4324 4438 4380
rect 4438 4324 4442 4380
rect 4378 4320 4442 4324
rect 4458 4380 4522 4384
rect 4458 4324 4462 4380
rect 4462 4324 4518 4380
rect 4518 4324 4522 4380
rect 4458 4320 4522 4324
rect 4538 4380 4602 4384
rect 4538 4324 4542 4380
rect 4542 4324 4598 4380
rect 4598 4324 4602 4380
rect 4538 4320 4602 4324
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 7805 4380 7869 4384
rect 7805 4324 7809 4380
rect 7809 4324 7865 4380
rect 7865 4324 7869 4380
rect 7805 4320 7869 4324
rect 7885 4380 7949 4384
rect 7885 4324 7889 4380
rect 7889 4324 7945 4380
rect 7945 4324 7949 4380
rect 7885 4320 7949 4324
rect 7965 4380 8029 4384
rect 7965 4324 7969 4380
rect 7969 4324 8025 4380
rect 8025 4324 8029 4380
rect 7965 4320 8029 4324
rect 8045 4380 8109 4384
rect 8045 4324 8049 4380
rect 8049 4324 8105 4380
rect 8105 4324 8109 4380
rect 8045 4320 8109 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 11392 4380 11456 4384
rect 11392 4324 11396 4380
rect 11396 4324 11452 4380
rect 11452 4324 11456 4380
rect 11392 4320 11456 4324
rect 11472 4380 11536 4384
rect 11472 4324 11476 4380
rect 11476 4324 11532 4380
rect 11532 4324 11536 4380
rect 11472 4320 11536 4324
rect 14659 4380 14723 4384
rect 14659 4324 14663 4380
rect 14663 4324 14719 4380
rect 14719 4324 14723 4380
rect 14659 4320 14723 4324
rect 14739 4380 14803 4384
rect 14739 4324 14743 4380
rect 14743 4324 14799 4380
rect 14799 4324 14803 4380
rect 14739 4320 14803 4324
rect 14819 4380 14883 4384
rect 14819 4324 14823 4380
rect 14823 4324 14879 4380
rect 14879 4324 14883 4380
rect 14819 4320 14883 4324
rect 14899 4380 14963 4384
rect 14899 4324 14903 4380
rect 14903 4324 14959 4380
rect 14959 4324 14963 4380
rect 14899 4320 14963 4324
rect 2665 3836 2729 3840
rect 2665 3780 2669 3836
rect 2669 3780 2725 3836
rect 2725 3780 2729 3836
rect 2665 3776 2729 3780
rect 2745 3836 2809 3840
rect 2745 3780 2749 3836
rect 2749 3780 2805 3836
rect 2805 3780 2809 3836
rect 2745 3776 2809 3780
rect 2825 3836 2889 3840
rect 2825 3780 2829 3836
rect 2829 3780 2885 3836
rect 2885 3780 2889 3836
rect 2825 3776 2889 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 9519 3836 9583 3840
rect 9519 3780 9523 3836
rect 9523 3780 9579 3836
rect 9579 3780 9583 3836
rect 9519 3776 9583 3780
rect 9599 3836 9663 3840
rect 9599 3780 9603 3836
rect 9603 3780 9659 3836
rect 9659 3780 9663 3836
rect 9599 3776 9663 3780
rect 9679 3836 9743 3840
rect 9679 3780 9683 3836
rect 9683 3780 9739 3836
rect 9739 3780 9743 3836
rect 9679 3776 9743 3780
rect 9759 3836 9823 3840
rect 9759 3780 9763 3836
rect 9763 3780 9819 3836
rect 9819 3780 9823 3836
rect 9759 3776 9823 3780
rect 12946 3836 13010 3840
rect 12946 3780 12950 3836
rect 12950 3780 13006 3836
rect 13006 3780 13010 3836
rect 12946 3776 13010 3780
rect 13026 3836 13090 3840
rect 13026 3780 13030 3836
rect 13030 3780 13086 3836
rect 13086 3780 13090 3836
rect 13026 3776 13090 3780
rect 13106 3836 13170 3840
rect 13106 3780 13110 3836
rect 13110 3780 13166 3836
rect 13166 3780 13170 3836
rect 13106 3776 13170 3780
rect 13186 3836 13250 3840
rect 13186 3780 13190 3836
rect 13190 3780 13246 3836
rect 13246 3780 13250 3836
rect 13186 3776 13250 3780
rect 4378 3292 4442 3296
rect 4378 3236 4382 3292
rect 4382 3236 4438 3292
rect 4438 3236 4442 3292
rect 4378 3232 4442 3236
rect 4458 3292 4522 3296
rect 4458 3236 4462 3292
rect 4462 3236 4518 3292
rect 4518 3236 4522 3292
rect 4458 3232 4522 3236
rect 4538 3292 4602 3296
rect 4538 3236 4542 3292
rect 4542 3236 4598 3292
rect 4598 3236 4602 3292
rect 4538 3232 4602 3236
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 7805 3292 7869 3296
rect 7805 3236 7809 3292
rect 7809 3236 7865 3292
rect 7865 3236 7869 3292
rect 7805 3232 7869 3236
rect 7885 3292 7949 3296
rect 7885 3236 7889 3292
rect 7889 3236 7945 3292
rect 7945 3236 7949 3292
rect 7885 3232 7949 3236
rect 7965 3292 8029 3296
rect 7965 3236 7969 3292
rect 7969 3236 8025 3292
rect 8025 3236 8029 3292
rect 7965 3232 8029 3236
rect 8045 3292 8109 3296
rect 8045 3236 8049 3292
rect 8049 3236 8105 3292
rect 8105 3236 8109 3292
rect 8045 3232 8109 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 11392 3292 11456 3296
rect 11392 3236 11396 3292
rect 11396 3236 11452 3292
rect 11452 3236 11456 3292
rect 11392 3232 11456 3236
rect 11472 3292 11536 3296
rect 11472 3236 11476 3292
rect 11476 3236 11532 3292
rect 11532 3236 11536 3292
rect 11472 3232 11536 3236
rect 14659 3292 14723 3296
rect 14659 3236 14663 3292
rect 14663 3236 14719 3292
rect 14719 3236 14723 3292
rect 14659 3232 14723 3236
rect 14739 3292 14803 3296
rect 14739 3236 14743 3292
rect 14743 3236 14799 3292
rect 14799 3236 14803 3292
rect 14739 3232 14803 3236
rect 14819 3292 14883 3296
rect 14819 3236 14823 3292
rect 14823 3236 14879 3292
rect 14879 3236 14883 3292
rect 14819 3232 14883 3236
rect 14899 3292 14963 3296
rect 14899 3236 14903 3292
rect 14903 3236 14959 3292
rect 14959 3236 14963 3292
rect 14899 3232 14963 3236
rect 2665 2748 2729 2752
rect 2665 2692 2669 2748
rect 2669 2692 2725 2748
rect 2725 2692 2729 2748
rect 2665 2688 2729 2692
rect 2745 2748 2809 2752
rect 2745 2692 2749 2748
rect 2749 2692 2805 2748
rect 2805 2692 2809 2748
rect 2745 2688 2809 2692
rect 2825 2748 2889 2752
rect 2825 2692 2829 2748
rect 2829 2692 2885 2748
rect 2885 2692 2889 2748
rect 2825 2688 2889 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 9519 2748 9583 2752
rect 9519 2692 9523 2748
rect 9523 2692 9579 2748
rect 9579 2692 9583 2748
rect 9519 2688 9583 2692
rect 9599 2748 9663 2752
rect 9599 2692 9603 2748
rect 9603 2692 9659 2748
rect 9659 2692 9663 2748
rect 9599 2688 9663 2692
rect 9679 2748 9743 2752
rect 9679 2692 9683 2748
rect 9683 2692 9739 2748
rect 9739 2692 9743 2748
rect 9679 2688 9743 2692
rect 9759 2748 9823 2752
rect 9759 2692 9763 2748
rect 9763 2692 9819 2748
rect 9819 2692 9823 2748
rect 9759 2688 9823 2692
rect 12946 2748 13010 2752
rect 12946 2692 12950 2748
rect 12950 2692 13006 2748
rect 13006 2692 13010 2748
rect 12946 2688 13010 2692
rect 13026 2748 13090 2752
rect 13026 2692 13030 2748
rect 13030 2692 13086 2748
rect 13086 2692 13090 2748
rect 13026 2688 13090 2692
rect 13106 2748 13170 2752
rect 13106 2692 13110 2748
rect 13110 2692 13166 2748
rect 13166 2692 13170 2748
rect 13106 2688 13170 2692
rect 13186 2748 13250 2752
rect 13186 2692 13190 2748
rect 13190 2692 13246 2748
rect 13246 2692 13250 2748
rect 13186 2688 13250 2692
rect 4378 2204 4442 2208
rect 4378 2148 4382 2204
rect 4382 2148 4438 2204
rect 4438 2148 4442 2204
rect 4378 2144 4442 2148
rect 4458 2204 4522 2208
rect 4458 2148 4462 2204
rect 4462 2148 4518 2204
rect 4518 2148 4522 2204
rect 4458 2144 4522 2148
rect 4538 2204 4602 2208
rect 4538 2148 4542 2204
rect 4542 2148 4598 2204
rect 4598 2148 4602 2204
rect 4538 2144 4602 2148
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 7805 2204 7869 2208
rect 7805 2148 7809 2204
rect 7809 2148 7865 2204
rect 7865 2148 7869 2204
rect 7805 2144 7869 2148
rect 7885 2204 7949 2208
rect 7885 2148 7889 2204
rect 7889 2148 7945 2204
rect 7945 2148 7949 2204
rect 7885 2144 7949 2148
rect 7965 2204 8029 2208
rect 7965 2148 7969 2204
rect 7969 2148 8025 2204
rect 8025 2148 8029 2204
rect 7965 2144 8029 2148
rect 8045 2204 8109 2208
rect 8045 2148 8049 2204
rect 8049 2148 8105 2204
rect 8105 2148 8109 2204
rect 8045 2144 8109 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 11392 2204 11456 2208
rect 11392 2148 11396 2204
rect 11396 2148 11452 2204
rect 11452 2148 11456 2204
rect 11392 2144 11456 2148
rect 11472 2204 11536 2208
rect 11472 2148 11476 2204
rect 11476 2148 11532 2204
rect 11532 2148 11536 2204
rect 11472 2144 11536 2148
rect 14659 2204 14723 2208
rect 14659 2148 14663 2204
rect 14663 2148 14719 2204
rect 14719 2148 14723 2204
rect 14659 2144 14723 2148
rect 14739 2204 14803 2208
rect 14739 2148 14743 2204
rect 14743 2148 14799 2204
rect 14799 2148 14803 2204
rect 14739 2144 14803 2148
rect 14819 2204 14883 2208
rect 14819 2148 14823 2204
rect 14823 2148 14879 2204
rect 14879 2148 14883 2204
rect 14819 2144 14883 2148
rect 14899 2204 14963 2208
rect 14899 2148 14903 2204
rect 14903 2148 14959 2204
rect 14959 2148 14963 2204
rect 14899 2144 14963 2148
<< metal4 >>
rect 2657 6016 2977 6576
rect 2657 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2977 6016
rect 2657 4928 2977 5952
rect 2657 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2977 4928
rect 2657 3840 2977 4864
rect 2657 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2977 3840
rect 2657 2752 2977 3776
rect 2657 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2977 2752
rect 2657 2128 2977 2688
rect 4370 6560 4690 6576
rect 4370 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4690 6560
rect 4370 5472 4690 6496
rect 4370 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4690 5472
rect 4370 4384 4690 5408
rect 4370 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4690 4384
rect 4370 3296 4690 4320
rect 4370 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4690 3296
rect 4370 2208 4690 3232
rect 4370 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4690 2208
rect 4370 2128 4690 2144
rect 6084 6016 6404 6576
rect 6084 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6404 6016
rect 6084 4928 6404 5952
rect 6084 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6404 4928
rect 6084 3840 6404 4864
rect 6084 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6404 3840
rect 6084 2752 6404 3776
rect 6084 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6404 2752
rect 6084 2128 6404 2688
rect 7797 6560 8117 6576
rect 7797 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8117 6560
rect 7797 5472 8117 6496
rect 7797 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8117 5472
rect 7797 4384 8117 5408
rect 7797 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8117 4384
rect 7797 3296 8117 4320
rect 7797 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8117 3296
rect 7797 2208 8117 3232
rect 7797 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8117 2208
rect 7797 2128 8117 2144
rect 9511 6016 9831 6576
rect 9511 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9831 6016
rect 9511 4928 9831 5952
rect 9511 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9831 4928
rect 9511 3840 9831 4864
rect 9511 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9831 3840
rect 9511 2752 9831 3776
rect 9511 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9831 2752
rect 9511 2128 9831 2688
rect 11224 6560 11544 6576
rect 11224 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11544 6560
rect 11224 5472 11544 6496
rect 11224 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11544 5472
rect 11224 4384 11544 5408
rect 11224 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11544 4384
rect 11224 3296 11544 4320
rect 11224 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11544 3296
rect 11224 2208 11544 3232
rect 11224 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11544 2208
rect 11224 2128 11544 2144
rect 12938 6016 13258 6576
rect 12938 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13258 6016
rect 12938 4928 13258 5952
rect 12938 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13258 4928
rect 12938 3840 13258 4864
rect 12938 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13258 3840
rect 12938 2752 13258 3776
rect 12938 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13258 2752
rect 12938 2128 13258 2688
rect 14651 6560 14971 6576
rect 14651 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14971 6560
rect 14651 5472 14971 6496
rect 14651 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14971 5472
rect 14651 4384 14971 5408
rect 14651 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14971 4384
rect 14651 3296 14971 4320
rect 14651 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14971 3296
rect 14651 2208 14971 3232
rect 14651 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14971 2208
rect 14651 2128 14971 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 1840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 2392 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 3680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 4232 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 4968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 1840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35
timestamp 1666464484
transform 1 0 4324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1666464484
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1666464484
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1666464484
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64
timestamp 1666464484
transform 1 0 6992 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp 1666464484
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1666464484
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1666464484
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94
timestamp 1666464484
transform 1 0 9752 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_102
timestamp 1666464484
transform 1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 1666464484
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_124
timestamp 1666464484
transform 1 0 12512 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_132
timestamp 1666464484
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1666464484
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1666464484
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1666464484
transform 1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7
timestamp 1666464484
transform 1 0 1748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19
timestamp 1666464484
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_73
timestamp 1666464484
transform 1 0 7820 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1666464484
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_8
timestamp 1666464484
transform 1 0 1840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_16
timestamp 1666464484
transform 1 0 2576 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1666464484
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1666464484
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1666464484
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_65
timestamp 1666464484
transform 1 0 7084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_70
timestamp 1666464484
transform 1 0 7544 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_77
timestamp 1666464484
transform 1 0 8188 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_84
timestamp 1666464484
transform 1 0 8832 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_96
timestamp 1666464484
transform 1 0 9936 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1666464484
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_145
timestamp 1666464484
transform 1 0 14444 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_8
timestamp 1666464484
transform 1 0 1840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1666464484
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_47
timestamp 1666464484
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_51
timestamp 1666464484
transform 1 0 5796 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_63
timestamp 1666464484
transform 1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_70
timestamp 1666464484
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1666464484
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_8
timestamp 1666464484
transform 1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_14
timestamp 1666464484
transform 1 0 2392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_18
timestamp 1666464484
transform 1 0 2760 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_21
timestamp 1666464484
transform 1 0 3036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_25
timestamp 1666464484
transform 1 0 3404 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1666464484
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_34
timestamp 1666464484
transform 1 0 4232 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_46
timestamp 1666464484
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1666464484
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_65
timestamp 1666464484
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_145
timestamp 1666464484
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1666464484
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_11
timestamp 1666464484
transform 1 0 2116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_18
timestamp 1666464484
transform 1 0 2760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_22
timestamp 1666464484
transform 1 0 3128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1666464484
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_36
timestamp 1666464484
transform 1 0 4416 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_42
timestamp 1666464484
transform 1 0 4968 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_54
timestamp 1666464484
transform 1 0 6072 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_66
timestamp 1666464484
transform 1 0 7176 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1666464484
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_145
timestamp 1666464484
transform 1 0 14444 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_12
timestamp 1666464484
transform 1 0 2208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1666464484
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_26
timestamp 1666464484
transform 1 0 3496 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_29
timestamp 1666464484
transform 1 0 3772 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_35
timestamp 1666464484
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_46
timestamp 1666464484
transform 1 0 5336 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1666464484
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_85
timestamp 1666464484
transform 1 0 8924 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_90
timestamp 1666464484
transform 1 0 9384 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_96
timestamp 1666464484
transform 1 0 9936 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1666464484
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_141
timestamp 1666464484
transform 1 0 14076 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_145
timestamp 1666464484
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_17
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_18
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_19
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1666464484
transform 1 0 3680 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1666464484
transform 1 0 8832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1666464484
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _00_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _01_
timestamp 1666464484
transform -1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _02_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp 1666464484
transform -1 0 4324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _04_
timestamp 1666464484
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp 1666464484
transform -1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1666464484
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp 1666464484
transform -1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1666464484
transform -1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1666464484
transform -1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1666464484
transform -1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform -1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform 1 0 9108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform -1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1666464484
transform -1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666464484
transform -1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1666464484
transform -1 0 3496 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1666464484
transform -1 0 3496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1666464484
transform -1 0 4416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1666464484
transform -1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666464484
transform -1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1666464484
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1666464484
transform 1 0 6624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1666464484
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1666464484
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1666464484
transform 1 0 10764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1666464484
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1666464484
transform 1 0 13432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1666464484
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1666464484
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 406 592
<< labels >>
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 ram_adrb[0]
port 0 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 ram_adrb[1]
port 1 nsew signal tristate
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 ram_adrb[2]
port 2 nsew signal tristate
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 ram_adrb[3]
port 3 nsew signal tristate
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 ram_adrb[4]
port 4 nsew signal tristate
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 ram_adrb[5]
port 5 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 ram_adrb[6]
port 6 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 ram_adrb[7]
port 7 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 ram_adrb[8]
port 8 nsew signal tristate
flabel metal2 s 1030 0 1086 800 0 FreeSans 224 90 0 0 ram_csb
port 9 nsew signal tristate
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 ram_web
port 10 nsew signal tristate
flabel metal4 s 2657 2128 2977 6576 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 6084 2128 6404 6576 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 9511 2128 9831 6576 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 12938 2128 13258 6576 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 4370 2128 4690 6576 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 7797 2128 8117 6576 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 11224 2128 11544 6576 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 14651 2128 14971 6576 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal2 s 386 8200 442 9000 0 FreeSans 224 90 0 0 wb_clk_i
port 13 nsew signal input
flabel metal2 s 1306 8200 1362 9000 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 14 nsew signal input
flabel metal2 s 5906 8200 5962 9000 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 15 nsew signal input
flabel metal2 s 6366 8200 6422 9000 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 16 nsew signal input
flabel metal2 s 6826 8200 6882 9000 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 17 nsew signal input
flabel metal2 s 7286 8200 7342 9000 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 18 nsew signal input
flabel metal2 s 7746 8200 7802 9000 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 19 nsew signal input
flabel metal2 s 8206 8200 8262 9000 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 20 nsew signal input
flabel metal2 s 8666 8200 8722 9000 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 21 nsew signal input
flabel metal2 s 9126 8200 9182 9000 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 22 nsew signal input
flabel metal2 s 9586 8200 9642 9000 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 23 nsew signal input
flabel metal2 s 10046 8200 10102 9000 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 24 nsew signal input
flabel metal2 s 1766 8200 1822 9000 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 25 nsew signal input
flabel metal2 s 10506 8200 10562 9000 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 26 nsew signal input
flabel metal2 s 10966 8200 11022 9000 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 27 nsew signal input
flabel metal2 s 11426 8200 11482 9000 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 28 nsew signal input
flabel metal2 s 11886 8200 11942 9000 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 29 nsew signal input
flabel metal2 s 12346 8200 12402 9000 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 30 nsew signal input
flabel metal2 s 12806 8200 12862 9000 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 31 nsew signal input
flabel metal2 s 13266 8200 13322 9000 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 32 nsew signal input
flabel metal2 s 13726 8200 13782 9000 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 33 nsew signal input
flabel metal2 s 14186 8200 14242 9000 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 34 nsew signal input
flabel metal2 s 14646 8200 14702 9000 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 35 nsew signal input
flabel metal2 s 2226 8200 2282 9000 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 36 nsew signal input
flabel metal2 s 15106 8200 15162 9000 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 37 nsew signal input
flabel metal2 s 15566 8200 15622 9000 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 38 nsew signal input
flabel metal2 s 2686 8200 2742 9000 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 39 nsew signal input
flabel metal2 s 3146 8200 3202 9000 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 40 nsew signal input
flabel metal2 s 3606 8200 3662 9000 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 41 nsew signal input
flabel metal2 s 4066 8200 4122 9000 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 42 nsew signal input
flabel metal2 s 4526 8200 4582 9000 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 43 nsew signal input
flabel metal2 s 4986 8200 5042 9000 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 44 nsew signal input
flabel metal2 s 5446 8200 5502 9000 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 45 nsew signal input
flabel metal2 s 846 8200 902 9000 0 FreeSans 224 90 0 0 wbs_we_i
port 46 nsew signal input
rlabel metal1 7958 5984 7958 5984 0 vccd1
rlabel via1 8037 6528 8037 6528 0 vssd1
rlabel metal1 2438 4114 2438 4114 0 net1
rlabel metal1 6716 3502 6716 3502 0 net10
rlabel metal2 2438 5066 2438 5066 0 net11
rlabel metal2 4002 3162 4002 3162 0 net12
rlabel metal2 5290 3162 5290 3162 0 net13
rlabel metal2 6670 3434 6670 3434 0 net14
rlabel metal1 7728 2414 7728 2414 0 net15
rlabel metal2 9430 3162 9430 3162 0 net16
rlabel metal2 10810 3434 10810 3434 0 net17
rlabel metal2 8694 3196 8694 3196 0 net18
rlabel metal2 7498 4352 7498 4352 0 net19
rlabel metal1 7544 4114 7544 4114 0 net2
rlabel metal2 14030 3196 14030 3196 0 net20
rlabel metal1 1886 2448 1886 2448 0 net21
rlabel metal2 2530 3434 2530 3434 0 net22
rlabel metal1 4094 4080 4094 4080 0 net3
rlabel metal1 4830 4590 4830 4590 0 net4
rlabel metal1 7038 5202 7038 5202 0 net5
rlabel metal2 8602 4964 8602 4964 0 net6
rlabel metal1 7958 4624 7958 4624 0 net7
rlabel metal1 7820 4114 7820 4114 0 net8
rlabel metal1 7038 4590 7038 4590 0 net9
rlabel metal2 3818 1520 3818 1520 0 ram_adrb[0]
rlabel metal2 5198 1520 5198 1520 0 ram_adrb[1]
rlabel metal2 6578 1520 6578 1520 0 ram_adrb[2]
rlabel metal2 7958 823 7958 823 0 ram_adrb[3]
rlabel metal2 9338 1520 9338 1520 0 ram_adrb[4]
rlabel metal2 10718 1520 10718 1520 0 ram_adrb[5]
rlabel metal2 12098 1520 12098 1520 0 ram_adrb[6]
rlabel metal2 13478 1520 13478 1520 0 ram_adrb[7]
rlabel metal2 14858 823 14858 823 0 ram_adrb[8]
rlabel metal2 1058 1520 1058 1520 0 ram_csb
rlabel metal2 2438 1520 2438 1520 0 ram_web
rlabel metal1 1472 5202 1472 5202 0 wbs_adr_i[0]
rlabel metal1 9016 6290 9016 6290 0 wbs_adr_i[16]
rlabel metal1 1840 5678 1840 5678 0 wbs_adr_i[1]
rlabel metal1 2116 6290 2116 6290 0 wbs_adr_i[2]
rlabel metal1 2668 6290 2668 6290 0 wbs_adr_i[3]
rlabel metal1 3220 5678 3220 5678 0 wbs_adr_i[4]
rlabel metal1 3450 6290 3450 6290 0 wbs_adr_i[5]
rlabel metal2 4186 6001 4186 6001 0 wbs_adr_i[6]
rlabel metal1 4600 6290 4600 6290 0 wbs_adr_i[7]
rlabel metal1 5060 6290 5060 6290 0 wbs_adr_i[8]
rlabel metal1 1288 4794 1288 4794 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 16000 9000
<< end >>
