// This is the unpowered netlist.
module tms1x00_ram (clk,
    wen,
    r_val,
    ram_addr,
    w_val);
 input clk;
 input wen;
 output [3:0] r_val;
 input [6:0] ram_addr;
 input [3:0] w_val;

 wire \RAM[0][0] ;
 wire \RAM[0][1] ;
 wire \RAM[0][2] ;
 wire \RAM[0][3] ;
 wire \RAM[100][0] ;
 wire \RAM[100][1] ;
 wire \RAM[100][2] ;
 wire \RAM[100][3] ;
 wire \RAM[101][0] ;
 wire \RAM[101][1] ;
 wire \RAM[101][2] ;
 wire \RAM[101][3] ;
 wire \RAM[102][0] ;
 wire \RAM[102][1] ;
 wire \RAM[102][2] ;
 wire \RAM[102][3] ;
 wire \RAM[103][0] ;
 wire \RAM[103][1] ;
 wire \RAM[103][2] ;
 wire \RAM[103][3] ;
 wire \RAM[104][0] ;
 wire \RAM[104][1] ;
 wire \RAM[104][2] ;
 wire \RAM[104][3] ;
 wire \RAM[105][0] ;
 wire \RAM[105][1] ;
 wire \RAM[105][2] ;
 wire \RAM[105][3] ;
 wire \RAM[106][0] ;
 wire \RAM[106][1] ;
 wire \RAM[106][2] ;
 wire \RAM[106][3] ;
 wire \RAM[107][0] ;
 wire \RAM[107][1] ;
 wire \RAM[107][2] ;
 wire \RAM[107][3] ;
 wire \RAM[108][0] ;
 wire \RAM[108][1] ;
 wire \RAM[108][2] ;
 wire \RAM[108][3] ;
 wire \RAM[109][0] ;
 wire \RAM[109][1] ;
 wire \RAM[109][2] ;
 wire \RAM[109][3] ;
 wire \RAM[10][0] ;
 wire \RAM[10][1] ;
 wire \RAM[10][2] ;
 wire \RAM[10][3] ;
 wire \RAM[110][0] ;
 wire \RAM[110][1] ;
 wire \RAM[110][2] ;
 wire \RAM[110][3] ;
 wire \RAM[111][0] ;
 wire \RAM[111][1] ;
 wire \RAM[111][2] ;
 wire \RAM[111][3] ;
 wire \RAM[112][0] ;
 wire \RAM[112][1] ;
 wire \RAM[112][2] ;
 wire \RAM[112][3] ;
 wire \RAM[113][0] ;
 wire \RAM[113][1] ;
 wire \RAM[113][2] ;
 wire \RAM[113][3] ;
 wire \RAM[114][0] ;
 wire \RAM[114][1] ;
 wire \RAM[114][2] ;
 wire \RAM[114][3] ;
 wire \RAM[115][0] ;
 wire \RAM[115][1] ;
 wire \RAM[115][2] ;
 wire \RAM[115][3] ;
 wire \RAM[116][0] ;
 wire \RAM[116][1] ;
 wire \RAM[116][2] ;
 wire \RAM[116][3] ;
 wire \RAM[117][0] ;
 wire \RAM[117][1] ;
 wire \RAM[117][2] ;
 wire \RAM[117][3] ;
 wire \RAM[118][0] ;
 wire \RAM[118][1] ;
 wire \RAM[118][2] ;
 wire \RAM[118][3] ;
 wire \RAM[119][0] ;
 wire \RAM[119][1] ;
 wire \RAM[119][2] ;
 wire \RAM[119][3] ;
 wire \RAM[11][0] ;
 wire \RAM[11][1] ;
 wire \RAM[11][2] ;
 wire \RAM[11][3] ;
 wire \RAM[120][0] ;
 wire \RAM[120][1] ;
 wire \RAM[120][2] ;
 wire \RAM[120][3] ;
 wire \RAM[121][0] ;
 wire \RAM[121][1] ;
 wire \RAM[121][2] ;
 wire \RAM[121][3] ;
 wire \RAM[122][0] ;
 wire \RAM[122][1] ;
 wire \RAM[122][2] ;
 wire \RAM[122][3] ;
 wire \RAM[123][0] ;
 wire \RAM[123][1] ;
 wire \RAM[123][2] ;
 wire \RAM[123][3] ;
 wire \RAM[124][0] ;
 wire \RAM[124][1] ;
 wire \RAM[124][2] ;
 wire \RAM[124][3] ;
 wire \RAM[125][0] ;
 wire \RAM[125][1] ;
 wire \RAM[125][2] ;
 wire \RAM[125][3] ;
 wire \RAM[126][0] ;
 wire \RAM[126][1] ;
 wire \RAM[126][2] ;
 wire \RAM[126][3] ;
 wire \RAM[127][0] ;
 wire \RAM[127][1] ;
 wire \RAM[127][2] ;
 wire \RAM[127][3] ;
 wire \RAM[12][0] ;
 wire \RAM[12][1] ;
 wire \RAM[12][2] ;
 wire \RAM[12][3] ;
 wire \RAM[13][0] ;
 wire \RAM[13][1] ;
 wire \RAM[13][2] ;
 wire \RAM[13][3] ;
 wire \RAM[14][0] ;
 wire \RAM[14][1] ;
 wire \RAM[14][2] ;
 wire \RAM[14][3] ;
 wire \RAM[15][0] ;
 wire \RAM[15][1] ;
 wire \RAM[15][2] ;
 wire \RAM[15][3] ;
 wire \RAM[16][0] ;
 wire \RAM[16][1] ;
 wire \RAM[16][2] ;
 wire \RAM[16][3] ;
 wire \RAM[17][0] ;
 wire \RAM[17][1] ;
 wire \RAM[17][2] ;
 wire \RAM[17][3] ;
 wire \RAM[18][0] ;
 wire \RAM[18][1] ;
 wire \RAM[18][2] ;
 wire \RAM[18][3] ;
 wire \RAM[19][0] ;
 wire \RAM[19][1] ;
 wire \RAM[19][2] ;
 wire \RAM[19][3] ;
 wire \RAM[1][0] ;
 wire \RAM[1][1] ;
 wire \RAM[1][2] ;
 wire \RAM[1][3] ;
 wire \RAM[20][0] ;
 wire \RAM[20][1] ;
 wire \RAM[20][2] ;
 wire \RAM[20][3] ;
 wire \RAM[21][0] ;
 wire \RAM[21][1] ;
 wire \RAM[21][2] ;
 wire \RAM[21][3] ;
 wire \RAM[22][0] ;
 wire \RAM[22][1] ;
 wire \RAM[22][2] ;
 wire \RAM[22][3] ;
 wire \RAM[23][0] ;
 wire \RAM[23][1] ;
 wire \RAM[23][2] ;
 wire \RAM[23][3] ;
 wire \RAM[24][0] ;
 wire \RAM[24][1] ;
 wire \RAM[24][2] ;
 wire \RAM[24][3] ;
 wire \RAM[25][0] ;
 wire \RAM[25][1] ;
 wire \RAM[25][2] ;
 wire \RAM[25][3] ;
 wire \RAM[26][0] ;
 wire \RAM[26][1] ;
 wire \RAM[26][2] ;
 wire \RAM[26][3] ;
 wire \RAM[27][0] ;
 wire \RAM[27][1] ;
 wire \RAM[27][2] ;
 wire \RAM[27][3] ;
 wire \RAM[28][0] ;
 wire \RAM[28][1] ;
 wire \RAM[28][2] ;
 wire \RAM[28][3] ;
 wire \RAM[29][0] ;
 wire \RAM[29][1] ;
 wire \RAM[29][2] ;
 wire \RAM[29][3] ;
 wire \RAM[2][0] ;
 wire \RAM[2][1] ;
 wire \RAM[2][2] ;
 wire \RAM[2][3] ;
 wire \RAM[30][0] ;
 wire \RAM[30][1] ;
 wire \RAM[30][2] ;
 wire \RAM[30][3] ;
 wire \RAM[31][0] ;
 wire \RAM[31][1] ;
 wire \RAM[31][2] ;
 wire \RAM[31][3] ;
 wire \RAM[32][0] ;
 wire \RAM[32][1] ;
 wire \RAM[32][2] ;
 wire \RAM[32][3] ;
 wire \RAM[33][0] ;
 wire \RAM[33][1] ;
 wire \RAM[33][2] ;
 wire \RAM[33][3] ;
 wire \RAM[34][0] ;
 wire \RAM[34][1] ;
 wire \RAM[34][2] ;
 wire \RAM[34][3] ;
 wire \RAM[35][0] ;
 wire \RAM[35][1] ;
 wire \RAM[35][2] ;
 wire \RAM[35][3] ;
 wire \RAM[36][0] ;
 wire \RAM[36][1] ;
 wire \RAM[36][2] ;
 wire \RAM[36][3] ;
 wire \RAM[37][0] ;
 wire \RAM[37][1] ;
 wire \RAM[37][2] ;
 wire \RAM[37][3] ;
 wire \RAM[38][0] ;
 wire \RAM[38][1] ;
 wire \RAM[38][2] ;
 wire \RAM[38][3] ;
 wire \RAM[39][0] ;
 wire \RAM[39][1] ;
 wire \RAM[39][2] ;
 wire \RAM[39][3] ;
 wire \RAM[3][0] ;
 wire \RAM[3][1] ;
 wire \RAM[3][2] ;
 wire \RAM[3][3] ;
 wire \RAM[40][0] ;
 wire \RAM[40][1] ;
 wire \RAM[40][2] ;
 wire \RAM[40][3] ;
 wire \RAM[41][0] ;
 wire \RAM[41][1] ;
 wire \RAM[41][2] ;
 wire \RAM[41][3] ;
 wire \RAM[42][0] ;
 wire \RAM[42][1] ;
 wire \RAM[42][2] ;
 wire \RAM[42][3] ;
 wire \RAM[43][0] ;
 wire \RAM[43][1] ;
 wire \RAM[43][2] ;
 wire \RAM[43][3] ;
 wire \RAM[44][0] ;
 wire \RAM[44][1] ;
 wire \RAM[44][2] ;
 wire \RAM[44][3] ;
 wire \RAM[45][0] ;
 wire \RAM[45][1] ;
 wire \RAM[45][2] ;
 wire \RAM[45][3] ;
 wire \RAM[46][0] ;
 wire \RAM[46][1] ;
 wire \RAM[46][2] ;
 wire \RAM[46][3] ;
 wire \RAM[47][0] ;
 wire \RAM[47][1] ;
 wire \RAM[47][2] ;
 wire \RAM[47][3] ;
 wire \RAM[48][0] ;
 wire \RAM[48][1] ;
 wire \RAM[48][2] ;
 wire \RAM[48][3] ;
 wire \RAM[49][0] ;
 wire \RAM[49][1] ;
 wire \RAM[49][2] ;
 wire \RAM[49][3] ;
 wire \RAM[4][0] ;
 wire \RAM[4][1] ;
 wire \RAM[4][2] ;
 wire \RAM[4][3] ;
 wire \RAM[50][0] ;
 wire \RAM[50][1] ;
 wire \RAM[50][2] ;
 wire \RAM[50][3] ;
 wire \RAM[51][0] ;
 wire \RAM[51][1] ;
 wire \RAM[51][2] ;
 wire \RAM[51][3] ;
 wire \RAM[52][0] ;
 wire \RAM[52][1] ;
 wire \RAM[52][2] ;
 wire \RAM[52][3] ;
 wire \RAM[53][0] ;
 wire \RAM[53][1] ;
 wire \RAM[53][2] ;
 wire \RAM[53][3] ;
 wire \RAM[54][0] ;
 wire \RAM[54][1] ;
 wire \RAM[54][2] ;
 wire \RAM[54][3] ;
 wire \RAM[55][0] ;
 wire \RAM[55][1] ;
 wire \RAM[55][2] ;
 wire \RAM[55][3] ;
 wire \RAM[56][0] ;
 wire \RAM[56][1] ;
 wire \RAM[56][2] ;
 wire \RAM[56][3] ;
 wire \RAM[57][0] ;
 wire \RAM[57][1] ;
 wire \RAM[57][2] ;
 wire \RAM[57][3] ;
 wire \RAM[58][0] ;
 wire \RAM[58][1] ;
 wire \RAM[58][2] ;
 wire \RAM[58][3] ;
 wire \RAM[59][0] ;
 wire \RAM[59][1] ;
 wire \RAM[59][2] ;
 wire \RAM[59][3] ;
 wire \RAM[5][0] ;
 wire \RAM[5][1] ;
 wire \RAM[5][2] ;
 wire \RAM[5][3] ;
 wire \RAM[60][0] ;
 wire \RAM[60][1] ;
 wire \RAM[60][2] ;
 wire \RAM[60][3] ;
 wire \RAM[61][0] ;
 wire \RAM[61][1] ;
 wire \RAM[61][2] ;
 wire \RAM[61][3] ;
 wire \RAM[62][0] ;
 wire \RAM[62][1] ;
 wire \RAM[62][2] ;
 wire \RAM[62][3] ;
 wire \RAM[63][0] ;
 wire \RAM[63][1] ;
 wire \RAM[63][2] ;
 wire \RAM[63][3] ;
 wire \RAM[64][0] ;
 wire \RAM[64][1] ;
 wire \RAM[64][2] ;
 wire \RAM[64][3] ;
 wire \RAM[65][0] ;
 wire \RAM[65][1] ;
 wire \RAM[65][2] ;
 wire \RAM[65][3] ;
 wire \RAM[66][0] ;
 wire \RAM[66][1] ;
 wire \RAM[66][2] ;
 wire \RAM[66][3] ;
 wire \RAM[67][0] ;
 wire \RAM[67][1] ;
 wire \RAM[67][2] ;
 wire \RAM[67][3] ;
 wire \RAM[68][0] ;
 wire \RAM[68][1] ;
 wire \RAM[68][2] ;
 wire \RAM[68][3] ;
 wire \RAM[69][0] ;
 wire \RAM[69][1] ;
 wire \RAM[69][2] ;
 wire \RAM[69][3] ;
 wire \RAM[6][0] ;
 wire \RAM[6][1] ;
 wire \RAM[6][2] ;
 wire \RAM[6][3] ;
 wire \RAM[70][0] ;
 wire \RAM[70][1] ;
 wire \RAM[70][2] ;
 wire \RAM[70][3] ;
 wire \RAM[71][0] ;
 wire \RAM[71][1] ;
 wire \RAM[71][2] ;
 wire \RAM[71][3] ;
 wire \RAM[72][0] ;
 wire \RAM[72][1] ;
 wire \RAM[72][2] ;
 wire \RAM[72][3] ;
 wire \RAM[73][0] ;
 wire \RAM[73][1] ;
 wire \RAM[73][2] ;
 wire \RAM[73][3] ;
 wire \RAM[74][0] ;
 wire \RAM[74][1] ;
 wire \RAM[74][2] ;
 wire \RAM[74][3] ;
 wire \RAM[75][0] ;
 wire \RAM[75][1] ;
 wire \RAM[75][2] ;
 wire \RAM[75][3] ;
 wire \RAM[76][0] ;
 wire \RAM[76][1] ;
 wire \RAM[76][2] ;
 wire \RAM[76][3] ;
 wire \RAM[77][0] ;
 wire \RAM[77][1] ;
 wire \RAM[77][2] ;
 wire \RAM[77][3] ;
 wire \RAM[78][0] ;
 wire \RAM[78][1] ;
 wire \RAM[78][2] ;
 wire \RAM[78][3] ;
 wire \RAM[79][0] ;
 wire \RAM[79][1] ;
 wire \RAM[79][2] ;
 wire \RAM[79][3] ;
 wire \RAM[7][0] ;
 wire \RAM[7][1] ;
 wire \RAM[7][2] ;
 wire \RAM[7][3] ;
 wire \RAM[80][0] ;
 wire \RAM[80][1] ;
 wire \RAM[80][2] ;
 wire \RAM[80][3] ;
 wire \RAM[81][0] ;
 wire \RAM[81][1] ;
 wire \RAM[81][2] ;
 wire \RAM[81][3] ;
 wire \RAM[82][0] ;
 wire \RAM[82][1] ;
 wire \RAM[82][2] ;
 wire \RAM[82][3] ;
 wire \RAM[83][0] ;
 wire \RAM[83][1] ;
 wire \RAM[83][2] ;
 wire \RAM[83][3] ;
 wire \RAM[84][0] ;
 wire \RAM[84][1] ;
 wire \RAM[84][2] ;
 wire \RAM[84][3] ;
 wire \RAM[85][0] ;
 wire \RAM[85][1] ;
 wire \RAM[85][2] ;
 wire \RAM[85][3] ;
 wire \RAM[86][0] ;
 wire \RAM[86][1] ;
 wire \RAM[86][2] ;
 wire \RAM[86][3] ;
 wire \RAM[87][0] ;
 wire \RAM[87][1] ;
 wire \RAM[87][2] ;
 wire \RAM[87][3] ;
 wire \RAM[88][0] ;
 wire \RAM[88][1] ;
 wire \RAM[88][2] ;
 wire \RAM[88][3] ;
 wire \RAM[89][0] ;
 wire \RAM[89][1] ;
 wire \RAM[89][2] ;
 wire \RAM[89][3] ;
 wire \RAM[8][0] ;
 wire \RAM[8][1] ;
 wire \RAM[8][2] ;
 wire \RAM[8][3] ;
 wire \RAM[90][0] ;
 wire \RAM[90][1] ;
 wire \RAM[90][2] ;
 wire \RAM[90][3] ;
 wire \RAM[91][0] ;
 wire \RAM[91][1] ;
 wire \RAM[91][2] ;
 wire \RAM[91][3] ;
 wire \RAM[92][0] ;
 wire \RAM[92][1] ;
 wire \RAM[92][2] ;
 wire \RAM[92][3] ;
 wire \RAM[93][0] ;
 wire \RAM[93][1] ;
 wire \RAM[93][2] ;
 wire \RAM[93][3] ;
 wire \RAM[94][0] ;
 wire \RAM[94][1] ;
 wire \RAM[94][2] ;
 wire \RAM[94][3] ;
 wire \RAM[95][0] ;
 wire \RAM[95][1] ;
 wire \RAM[95][2] ;
 wire \RAM[95][3] ;
 wire \RAM[96][0] ;
 wire \RAM[96][1] ;
 wire \RAM[96][2] ;
 wire \RAM[96][3] ;
 wire \RAM[97][0] ;
 wire \RAM[97][1] ;
 wire \RAM[97][2] ;
 wire \RAM[97][3] ;
 wire \RAM[98][0] ;
 wire \RAM[98][1] ;
 wire \RAM[98][2] ;
 wire \RAM[98][3] ;
 wire \RAM[99][0] ;
 wire \RAM[99][1] ;
 wire \RAM[99][2] ;
 wire \RAM[99][3] ;
 wire \RAM[9][0] ;
 wire \RAM[9][1] ;
 wire \RAM[9][2] ;
 wire \RAM[9][3] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__or2_1 _1628_ (.A(net5),
    .B(net6),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_4 _1629_ (.A(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_4 _1630_ (.A(net4),
    .X(_0514_));
 sky130_fd_sc_hd__buf_2 _1631_ (.A(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__buf_4 _1632_ (.A(net2),
    .X(_0516_));
 sky130_fd_sc_hd__buf_4 _1633_ (.A(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_4 _1634_ (.A(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__buf_6 _1635_ (.A(net1),
    .X(_0519_));
 sky130_fd_sc_hd__buf_6 _1636_ (.A(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__buf_6 _1637_ (.A(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _1638_ (.A0(\RAM[70][0] ),
    .A1(\RAM[71][0] ),
    .S(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__clkinv_2 _1639_ (.A(net2),
    .Y(_0523_));
 sky130_fd_sc_hd__clkbuf_4 _1640_ (.A(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__buf_2 _1641_ (.A(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__clkbuf_8 _1642_ (.A(net1),
    .X(_0526_));
 sky130_fd_sc_hd__buf_6 _1643_ (.A(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_8 _1644_ (.A(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _1645_ (.A0(\RAM[68][0] ),
    .A1(\RAM[69][0] ),
    .S(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__inv_2 _1646_ (.A(net3),
    .Y(_0530_));
 sky130_fd_sc_hd__clkbuf_4 _1647_ (.A(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__a21o_1 _1648_ (.A1(_0525_),
    .A2(_0529_),
    .B1(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__a21oi_1 _1649_ (.A1(_0518_),
    .A2(_0522_),
    .B1(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__buf_2 _1650_ (.A(net3),
    .X(_0534_));
 sky130_fd_sc_hd__clkbuf_4 _1651_ (.A(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__buf_2 _1652_ (.A(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__buf_6 _1653_ (.A(net1),
    .X(_0537_));
 sky130_fd_sc_hd__buf_8 _1654_ (.A(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__buf_4 _1655_ (.A(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__mux4_1 _1656_ (.A0(\RAM[64][0] ),
    .A1(\RAM[65][0] ),
    .A2(\RAM[66][0] ),
    .A3(\RAM[67][0] ),
    .S0(_0539_),
    .S1(_0517_),
    .X(_0540_));
 sky130_fd_sc_hd__nor2_1 _1657_ (.A(_0536_),
    .B(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__mux2_1 _1658_ (.A0(\RAM[78][0] ),
    .A1(\RAM[79][0] ),
    .S(_0521_),
    .X(_0542_));
 sky130_fd_sc_hd__buf_6 _1659_ (.A(_0526_),
    .X(_0543_));
 sky130_fd_sc_hd__buf_6 _1660_ (.A(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _1661_ (.A0(\RAM[76][0] ),
    .A1(\RAM[77][0] ),
    .S(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__a21o_1 _1662_ (.A1(_0525_),
    .A2(_0545_),
    .B1(_0531_),
    .X(_0546_));
 sky130_fd_sc_hd__a21oi_1 _1663_ (.A1(_0518_),
    .A2(_0542_),
    .B1(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__clkbuf_8 _1664_ (.A(net2),
    .X(_0548_));
 sky130_fd_sc_hd__buf_6 _1665_ (.A(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__buf_4 _1666_ (.A(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__mux4_1 _1667_ (.A0(\RAM[72][0] ),
    .A1(\RAM[73][0] ),
    .A2(\RAM[74][0] ),
    .A3(\RAM[75][0] ),
    .S0(_0539_),
    .S1(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__o21ai_1 _1668_ (.A1(_0536_),
    .A2(_0551_),
    .B1(_0515_),
    .Y(_0552_));
 sky130_fd_sc_hd__o32a_1 _1669_ (.A1(_0515_),
    .A2(_0533_),
    .A3(_0541_),
    .B1(_0547_),
    .B2(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__nor2_1 _1670_ (.A(_0513_),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__inv_2 _1671_ (.A(net7),
    .Y(_0555_));
 sky130_fd_sc_hd__or2_1 _1672_ (.A(_0534_),
    .B(net4),
    .X(_0556_));
 sky130_fd_sc_hd__clkbuf_4 _1673_ (.A(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__buf_4 _1674_ (.A(_0548_),
    .X(_0558_));
 sky130_fd_sc_hd__mux4_1 _1675_ (.A0(\RAM[112][0] ),
    .A1(\RAM[113][0] ),
    .A2(\RAM[114][0] ),
    .A3(\RAM[115][0] ),
    .S0(_0528_),
    .S1(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__or2b_1 _1676_ (.A(_0534_),
    .B_N(_0514_),
    .X(_0560_));
 sky130_fd_sc_hd__buf_4 _1677_ (.A(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__mux4_1 _1678_ (.A0(\RAM[120][0] ),
    .A1(\RAM[121][0] ),
    .A2(\RAM[122][0] ),
    .A3(\RAM[123][0] ),
    .S0(_0527_),
    .S1(_0548_),
    .X(_0562_));
 sky130_fd_sc_hd__nand2_1 _1679_ (.A(_0534_),
    .B(_0514_),
    .Y(_0563_));
 sky130_fd_sc_hd__buf_6 _1680_ (.A(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__buf_6 _1681_ (.A(_0526_),
    .X(_0565_));
 sky130_fd_sc_hd__buf_4 _1682_ (.A(net2),
    .X(_0566_));
 sky130_fd_sc_hd__mux4_1 _1683_ (.A0(\RAM[124][0] ),
    .A1(\RAM[125][0] ),
    .A2(\RAM[126][0] ),
    .A3(\RAM[127][0] ),
    .S0(_0565_),
    .S1(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__o22a_1 _1684_ (.A1(_0561_),
    .A2(_0562_),
    .B1(_0564_),
    .B2(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__or2b_1 _1685_ (.A(net4),
    .B_N(_0534_),
    .X(_0569_));
 sky130_fd_sc_hd__buf_4 _1686_ (.A(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__buf_6 _1687_ (.A(_0526_),
    .X(_0571_));
 sky130_fd_sc_hd__mux4_1 _1688_ (.A0(\RAM[116][0] ),
    .A1(\RAM[117][0] ),
    .A2(\RAM[118][0] ),
    .A3(\RAM[119][0] ),
    .S0(_0571_),
    .S1(_0516_),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_4 _1689_ (.A(net5),
    .X(_0573_));
 sky130_fd_sc_hd__nand2_4 _1690_ (.A(_0573_),
    .B(net6),
    .Y(_0574_));
 sky130_fd_sc_hd__o21ba_1 _1691_ (.A1(_0570_),
    .A2(_0572_),
    .B1_N(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__o211a_1 _1692_ (.A1(_0557_),
    .A2(_0559_),
    .B1(_0568_),
    .C1(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__and2_1 _1693_ (.A(_0530_),
    .B(_0514_),
    .X(_0577_));
 sky130_fd_sc_hd__buf_4 _1694_ (.A(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _1695_ (.A0(\RAM[104][0] ),
    .A1(\RAM[105][0] ),
    .S(_0526_),
    .X(_0579_));
 sky130_fd_sc_hd__or2_1 _1696_ (.A(_0516_),
    .B(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _1697_ (.A0(\RAM[106][0] ),
    .A1(\RAM[107][0] ),
    .S(_0537_),
    .X(_0581_));
 sky130_fd_sc_hd__or2_1 _1698_ (.A(_0523_),
    .B(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__mux4_1 _1699_ (.A0(\RAM[96][0] ),
    .A1(\RAM[97][0] ),
    .A2(\RAM[98][0] ),
    .A3(\RAM[99][0] ),
    .S0(_0565_),
    .S1(_0516_),
    .X(_0583_));
 sky130_fd_sc_hd__nor2_4 _1700_ (.A(_0534_),
    .B(_0514_),
    .Y(_0584_));
 sky130_fd_sc_hd__a32o_1 _1701_ (.A1(_0578_),
    .A2(_0580_),
    .A3(_0582_),
    .B1(_0583_),
    .B2(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__and2_1 _1702_ (.A(_0534_),
    .B(_0514_),
    .X(_0586_));
 sky130_fd_sc_hd__clkbuf_4 _1703_ (.A(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__mux4_1 _1704_ (.A0(\RAM[108][0] ),
    .A1(\RAM[109][0] ),
    .A2(\RAM[110][0] ),
    .A3(\RAM[111][0] ),
    .S0(_0527_),
    .S1(_0566_),
    .X(_0588_));
 sky130_fd_sc_hd__mux4_1 _1705_ (.A0(\RAM[100][0] ),
    .A1(\RAM[101][0] ),
    .A2(\RAM[102][0] ),
    .A3(\RAM[103][0] ),
    .S0(_0571_),
    .S1(_0516_),
    .X(_0589_));
 sky130_fd_sc_hd__and2b_2 _1706_ (.A_N(_0514_),
    .B(_0534_),
    .X(_0590_));
 sky130_fd_sc_hd__a22o_1 _1707_ (.A1(_0587_),
    .A2(_0588_),
    .B1(_0589_),
    .B2(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__and2b_1 _1708_ (.A_N(_0573_),
    .B(net6),
    .X(_0592_));
 sky130_fd_sc_hd__o21a_1 _1709_ (.A1(_0585_),
    .A2(_0591_),
    .B1(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__mux4_1 _1710_ (.A0(\RAM[84][0] ),
    .A1(\RAM[85][0] ),
    .A2(\RAM[86][0] ),
    .A3(\RAM[87][0] ),
    .S0(_0565_),
    .S1(_0566_),
    .X(_0594_));
 sky130_fd_sc_hd__buf_4 _1711_ (.A(net2),
    .X(_0595_));
 sky130_fd_sc_hd__mux4_1 _1712_ (.A0(\RAM[88][0] ),
    .A1(\RAM[89][0] ),
    .A2(\RAM[90][0] ),
    .A3(\RAM[91][0] ),
    .S0(_0543_),
    .S1(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__a22o_1 _1713_ (.A1(_0590_),
    .A2(_0594_),
    .B1(_0596_),
    .B2(_0578_),
    .X(_0597_));
 sky130_fd_sc_hd__mux4_1 _1714_ (.A0(\RAM[92][0] ),
    .A1(\RAM[93][0] ),
    .A2(\RAM[94][0] ),
    .A3(\RAM[95][0] ),
    .S0(_0565_),
    .S1(_0516_),
    .X(_0598_));
 sky130_fd_sc_hd__mux4_1 _1715_ (.A0(\RAM[80][0] ),
    .A1(\RAM[81][0] ),
    .A2(\RAM[82][0] ),
    .A3(\RAM[83][0] ),
    .S0(_0543_),
    .S1(_0595_),
    .X(_0599_));
 sky130_fd_sc_hd__a22o_1 _1716_ (.A1(_0587_),
    .A2(_0598_),
    .B1(_0599_),
    .B2(_0584_),
    .X(_0600_));
 sky130_fd_sc_hd__or2b_1 _1717_ (.A(net6),
    .B_N(_0573_),
    .X(_0601_));
 sky130_fd_sc_hd__buf_2 _1718_ (.A(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__o21ba_1 _1719_ (.A1(_0597_),
    .A2(_0600_),
    .B1_N(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__or4_1 _1720_ (.A(_0555_),
    .B(_0576_),
    .C(_0593_),
    .D(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__nor2_1 _1721_ (.A(_0573_),
    .B(net6),
    .Y(_0605_));
 sky130_fd_sc_hd__buf_6 _1722_ (.A(_0526_),
    .X(_0606_));
 sky130_fd_sc_hd__buf_4 _1723_ (.A(net2),
    .X(_0607_));
 sky130_fd_sc_hd__buf_4 _1724_ (.A(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__mux4_1 _1725_ (.A0(\RAM[8][0] ),
    .A1(\RAM[9][0] ),
    .A2(\RAM[10][0] ),
    .A3(\RAM[11][0] ),
    .S0(_0606_),
    .S1(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__or2_1 _1726_ (.A(_0535_),
    .B(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__buf_4 _1727_ (.A(_0565_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _1728_ (.A0(\RAM[14][0] ),
    .A1(\RAM[15][0] ),
    .S(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _1729_ (.A0(\RAM[12][0] ),
    .A1(\RAM[13][0] ),
    .S(_0571_),
    .X(_0613_));
 sky130_fd_sc_hd__buf_4 _1730_ (.A(_0530_),
    .X(_0614_));
 sky130_fd_sc_hd__a21o_1 _1731_ (.A1(_0524_),
    .A2(_0613_),
    .B1(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__a21o_1 _1732_ (.A1(_0550_),
    .A2(_0612_),
    .B1(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _1733_ (.A0(\RAM[4][0] ),
    .A1(\RAM[5][0] ),
    .S(_0528_),
    .X(_0617_));
 sky130_fd_sc_hd__buf_6 _1734_ (.A(_0548_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _1735_ (.A0(\RAM[6][0] ),
    .A1(\RAM[7][0] ),
    .S(_0527_),
    .X(_0619_));
 sky130_fd_sc_hd__and2_1 _1736_ (.A(_0618_),
    .B(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__a211o_1 _1737_ (.A1(_0525_),
    .A2(_0617_),
    .B1(_0620_),
    .C1(_0531_),
    .X(_0621_));
 sky130_fd_sc_hd__buf_8 _1738_ (.A(_0537_),
    .X(_0622_));
 sky130_fd_sc_hd__mux4_1 _1739_ (.A0(\RAM[0][0] ),
    .A1(\RAM[1][0] ),
    .A2(\RAM[2][0] ),
    .A3(\RAM[3][0] ),
    .S0(_0622_),
    .S1(_0549_),
    .X(_0623_));
 sky130_fd_sc_hd__clkbuf_4 _1740_ (.A(_0514_),
    .X(_0624_));
 sky130_fd_sc_hd__o21ba_1 _1741_ (.A1(_0535_),
    .A2(_0623_),
    .B1_N(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__a32o_1 _1742_ (.A1(_0515_),
    .A2(_0610_),
    .A3(_0616_),
    .B1(_0621_),
    .B2(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__buf_4 _1743_ (.A(_0590_),
    .X(_0627_));
 sky130_fd_sc_hd__buf_8 _1744_ (.A(_0607_),
    .X(_0628_));
 sky130_fd_sc_hd__mux4_1 _1745_ (.A0(\RAM[20][0] ),
    .A1(\RAM[21][0] ),
    .A2(\RAM[22][0] ),
    .A3(\RAM[23][0] ),
    .S0(_0538_),
    .S1(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__mux4_1 _1746_ (.A0(\RAM[24][0] ),
    .A1(\RAM[25][0] ),
    .A2(\RAM[26][0] ),
    .A3(\RAM[27][0] ),
    .S0(_0622_),
    .S1(_0549_),
    .X(_0630_));
 sky130_fd_sc_hd__a22o_1 _1747_ (.A1(_0627_),
    .A2(_0629_),
    .B1(_0630_),
    .B2(_0578_),
    .X(_0631_));
 sky130_fd_sc_hd__mux4_1 _1748_ (.A0(\RAM[28][0] ),
    .A1(\RAM[29][0] ),
    .A2(\RAM[30][0] ),
    .A3(\RAM[31][0] ),
    .S0(_0538_),
    .S1(_0628_),
    .X(_0632_));
 sky130_fd_sc_hd__mux4_1 _1749_ (.A0(\RAM[16][0] ),
    .A1(\RAM[17][0] ),
    .A2(\RAM[18][0] ),
    .A3(\RAM[19][0] ),
    .S0(_0622_),
    .S1(_0549_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_4 _1750_ (.A(_0584_),
    .X(_0634_));
 sky130_fd_sc_hd__a22o_1 _1751_ (.A1(_0587_),
    .A2(_0632_),
    .B1(_0633_),
    .B2(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__o21ba_1 _1752_ (.A1(_0631_),
    .A2(_0635_),
    .B1_N(_0602_),
    .X(_0636_));
 sky130_fd_sc_hd__buf_8 _1753_ (.A(_0526_),
    .X(_0637_));
 sky130_fd_sc_hd__buf_6 _1754_ (.A(_0607_),
    .X(_0638_));
 sky130_fd_sc_hd__mux4_1 _1755_ (.A0(\RAM[44][0] ),
    .A1(\RAM[45][0] ),
    .A2(\RAM[46][0] ),
    .A3(\RAM[47][0] ),
    .S0(_0637_),
    .S1(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__mux4_1 _1756_ (.A0(\RAM[40][0] ),
    .A1(\RAM[41][0] ),
    .A2(\RAM[42][0] ),
    .A3(\RAM[43][0] ),
    .S0(_0526_),
    .S1(net2),
    .X(_0640_));
 sky130_fd_sc_hd__or2_1 _1757_ (.A(_0535_),
    .B(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__o211a_1 _1758_ (.A1(_0531_),
    .A2(_0639_),
    .B1(_0641_),
    .C1(_0624_),
    .X(_0642_));
 sky130_fd_sc_hd__mux4_1 _1759_ (.A0(\RAM[32][0] ),
    .A1(\RAM[33][0] ),
    .A2(\RAM[34][0] ),
    .A3(\RAM[35][0] ),
    .S0(_0606_),
    .S1(_0608_),
    .X(_0643_));
 sky130_fd_sc_hd__mux4_1 _1760_ (.A0(\RAM[36][0] ),
    .A1(\RAM[37][0] ),
    .A2(\RAM[38][0] ),
    .A3(\RAM[39][0] ),
    .S0(_0538_),
    .S1(_0628_),
    .X(_0644_));
 sky130_fd_sc_hd__a22o_1 _1761_ (.A1(_0634_),
    .A2(_0643_),
    .B1(_0644_),
    .B2(_0627_),
    .X(_0645_));
 sky130_fd_sc_hd__mux4_1 _1762_ (.A0(\RAM[52][0] ),
    .A1(\RAM[53][0] ),
    .A2(\RAM[54][0] ),
    .A3(\RAM[55][0] ),
    .S0(_0537_),
    .S1(_0607_),
    .X(_0646_));
 sky130_fd_sc_hd__mux4_1 _1763_ (.A0(\RAM[56][0] ),
    .A1(\RAM[57][0] ),
    .A2(\RAM[58][0] ),
    .A3(\RAM[59][0] ),
    .S0(_0519_),
    .S1(_0548_),
    .X(_0647_));
 sky130_fd_sc_hd__o22a_1 _1764_ (.A1(_0570_),
    .A2(_0646_),
    .B1(_0647_),
    .B2(_0561_),
    .X(_0648_));
 sky130_fd_sc_hd__mux4_1 _1765_ (.A0(\RAM[60][0] ),
    .A1(\RAM[61][0] ),
    .A2(\RAM[62][0] ),
    .A3(\RAM[63][0] ),
    .S0(_0537_),
    .S1(_0607_),
    .X(_0649_));
 sky130_fd_sc_hd__mux4_1 _1766_ (.A0(\RAM[48][0] ),
    .A1(\RAM[49][0] ),
    .A2(\RAM[50][0] ),
    .A3(\RAM[51][0] ),
    .S0(_0519_),
    .S1(_0607_),
    .X(_0650_));
 sky130_fd_sc_hd__o22a_1 _1767_ (.A1(_0564_),
    .A2(_0649_),
    .B1(_0650_),
    .B2(_0557_),
    .X(_0651_));
 sky130_fd_sc_hd__a21bo_1 _1768_ (.A1(_0648_),
    .A2(_0651_),
    .B1_N(_0573_),
    .X(_0652_));
 sky130_fd_sc_hd__o311a_1 _1769_ (.A1(_0573_),
    .A2(_0642_),
    .A3(_0645_),
    .B1(_0652_),
    .C1(net6),
    .X(_0653_));
 sky130_fd_sc_hd__a211o_1 _1770_ (.A1(_0605_),
    .A2(_0626_),
    .B1(_0636_),
    .C1(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__o22a_1 _1771_ (.A1(_0554_),
    .A2(_0604_),
    .B1(_0654_),
    .B2(net7),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 _1772_ (.A0(\RAM[60][1] ),
    .A1(\RAM[61][1] ),
    .A2(\RAM[62][1] ),
    .A3(\RAM[63][1] ),
    .S0(_0521_),
    .S1(_0550_),
    .X(_0655_));
 sky130_fd_sc_hd__mux4_1 _1773_ (.A0(\RAM[48][1] ),
    .A1(\RAM[49][1] ),
    .A2(\RAM[50][1] ),
    .A3(\RAM[51][1] ),
    .S0(_0521_),
    .S1(_0550_),
    .X(_0656_));
 sky130_fd_sc_hd__mux4_1 _1774_ (.A0(\RAM[52][1] ),
    .A1(\RAM[53][1] ),
    .A2(\RAM[54][1] ),
    .A3(\RAM[55][1] ),
    .S0(_0520_),
    .S1(_0618_),
    .X(_0657_));
 sky130_fd_sc_hd__mux4_1 _1775_ (.A0(\RAM[56][1] ),
    .A1(\RAM[57][1] ),
    .A2(\RAM[58][1] ),
    .A3(\RAM[59][1] ),
    .S0(_0528_),
    .S1(_0558_),
    .X(_0658_));
 sky130_fd_sc_hd__o22a_1 _1776_ (.A1(_0570_),
    .A2(_0657_),
    .B1(_0658_),
    .B2(_0561_),
    .X(_0659_));
 sky130_fd_sc_hd__o221ai_2 _1777_ (.A1(_0564_),
    .A2(_0655_),
    .B1(_0656_),
    .B2(_0557_),
    .C1(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__mux4_1 _1778_ (.A0(\RAM[36][1] ),
    .A1(\RAM[37][1] ),
    .A2(\RAM[38][1] ),
    .A3(\RAM[39][1] ),
    .S0(_0538_),
    .S1(_0628_),
    .X(_0661_));
 sky130_fd_sc_hd__mux4_1 _1779_ (.A0(\RAM[32][1] ),
    .A1(\RAM[33][1] ),
    .A2(\RAM[34][1] ),
    .A3(\RAM[35][1] ),
    .S0(_0606_),
    .S1(_0608_),
    .X(_0662_));
 sky130_fd_sc_hd__mux4_1 _1780_ (.A0(\RAM[44][1] ),
    .A1(\RAM[45][1] ),
    .A2(\RAM[46][1] ),
    .A3(\RAM[47][1] ),
    .S0(_0606_),
    .S1(_0628_),
    .X(_0663_));
 sky130_fd_sc_hd__mux4_1 _1781_ (.A0(\RAM[40][1] ),
    .A1(\RAM[41][1] ),
    .A2(\RAM[42][1] ),
    .A3(\RAM[43][1] ),
    .S0(_0538_),
    .S1(_0628_),
    .X(_0664_));
 sky130_fd_sc_hd__mux4_1 _1782_ (.A0(_0661_),
    .A1(_0662_),
    .A2(_0663_),
    .A3(_0664_),
    .S0(_0614_),
    .S1(_0624_),
    .X(_0665_));
 sky130_fd_sc_hd__o21ai_1 _1783_ (.A1(_0573_),
    .A2(_0665_),
    .B1(net6),
    .Y(_0666_));
 sky130_fd_sc_hd__a21o_1 _1784_ (.A1(_0573_),
    .A2(_0660_),
    .B1(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__mux4_1 _1785_ (.A0(\RAM[0][1] ),
    .A1(\RAM[1][1] ),
    .A2(\RAM[2][1] ),
    .A3(\RAM[3][1] ),
    .S0(_0565_),
    .S1(_0566_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _1786_ (.A0(\RAM[6][1] ),
    .A1(\RAM[7][1] ),
    .S(_0565_),
    .X(_0669_));
 sky130_fd_sc_hd__nand2_1 _1787_ (.A(_0558_),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__mux2_1 _1788_ (.A0(\RAM[4][1] ),
    .A1(\RAM[5][1] ),
    .S(_0519_),
    .X(_0671_));
 sky130_fd_sc_hd__a21oi_1 _1789_ (.A1(_0524_),
    .A2(_0671_),
    .B1(_0530_),
    .Y(_0672_));
 sky130_fd_sc_hd__a2bb2o_1 _1790_ (.A1_N(_0535_),
    .A2_N(_0668_),
    .B1(_0670_),
    .B2(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _1791_ (.A0(\RAM[14][1] ),
    .A1(\RAM[15][1] ),
    .S(_0611_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _1792_ (.A0(\RAM[12][1] ),
    .A1(\RAM[13][1] ),
    .S(_0637_),
    .X(_0675_));
 sky130_fd_sc_hd__a21o_1 _1793_ (.A1(_0524_),
    .A2(_0675_),
    .B1(_0614_),
    .X(_0676_));
 sky130_fd_sc_hd__a21oi_1 _1794_ (.A1(_0518_),
    .A2(_0674_),
    .B1(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__mux4_1 _1795_ (.A0(\RAM[8][1] ),
    .A1(\RAM[9][1] ),
    .A2(\RAM[10][1] ),
    .A3(\RAM[11][1] ),
    .S0(_0622_),
    .S1(_0549_),
    .X(_0678_));
 sky130_fd_sc_hd__o21ai_1 _1796_ (.A1(_0536_),
    .A2(_0678_),
    .B1(_0624_),
    .Y(_0679_));
 sky130_fd_sc_hd__o22a_1 _1797_ (.A1(_0624_),
    .A2(_0673_),
    .B1(_0677_),
    .B2(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__mux4_1 _1798_ (.A0(\RAM[20][1] ),
    .A1(\RAM[21][1] ),
    .A2(\RAM[22][1] ),
    .A3(\RAM[23][1] ),
    .S0(_0622_),
    .S1(_0549_),
    .X(_0681_));
 sky130_fd_sc_hd__mux4_1 _1799_ (.A0(\RAM[24][1] ),
    .A1(\RAM[25][1] ),
    .A2(\RAM[26][1] ),
    .A3(\RAM[27][1] ),
    .S0(_0520_),
    .S1(_0618_),
    .X(_0682_));
 sky130_fd_sc_hd__a22o_1 _1800_ (.A1(_0627_),
    .A2(_0681_),
    .B1(_0682_),
    .B2(_0578_),
    .X(_0683_));
 sky130_fd_sc_hd__mux4_1 _1801_ (.A0(\RAM[28][1] ),
    .A1(\RAM[29][1] ),
    .A2(\RAM[30][1] ),
    .A3(\RAM[31][1] ),
    .S0(_0520_),
    .S1(_0618_),
    .X(_0684_));
 sky130_fd_sc_hd__mux4_1 _1802_ (.A0(\RAM[16][1] ),
    .A1(\RAM[17][1] ),
    .A2(\RAM[18][1] ),
    .A3(\RAM[19][1] ),
    .S0(_0520_),
    .S1(_0618_),
    .X(_0685_));
 sky130_fd_sc_hd__a22o_1 _1803_ (.A1(_0587_),
    .A2(_0684_),
    .B1(_0685_),
    .B2(_0634_),
    .X(_0686_));
 sky130_fd_sc_hd__nor2_1 _1804_ (.A(_0683_),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__o221a_1 _1805_ (.A1(_0513_),
    .A2(_0680_),
    .B1(_0687_),
    .B2(_0602_),
    .C1(_0555_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _1806_ (.A0(\RAM[70][1] ),
    .A1(\RAM[71][1] ),
    .S(_0520_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _1807_ (.A0(\RAM[68][1] ),
    .A1(\RAM[69][1] ),
    .S(_0565_),
    .X(_0690_));
 sky130_fd_sc_hd__a21o_1 _1808_ (.A1(_0524_),
    .A2(_0690_),
    .B1(_0530_),
    .X(_0691_));
 sky130_fd_sc_hd__a21oi_1 _1809_ (.A1(_0550_),
    .A2(_0689_),
    .B1(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__mux4_1 _1810_ (.A0(\RAM[64][1] ),
    .A1(\RAM[65][1] ),
    .A2(\RAM[66][1] ),
    .A3(\RAM[67][1] ),
    .S0(_0622_),
    .S1(_0549_),
    .X(_0693_));
 sky130_fd_sc_hd__nor2_1 _1811_ (.A(_0535_),
    .B(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__mux2_1 _1812_ (.A0(\RAM[78][1] ),
    .A1(\RAM[79][1] ),
    .S(_0544_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _1813_ (.A0(\RAM[76][1] ),
    .A1(\RAM[77][1] ),
    .S(_0606_),
    .X(_0696_));
 sky130_fd_sc_hd__a21o_1 _1814_ (.A1(_0525_),
    .A2(_0696_),
    .B1(_0614_),
    .X(_0697_));
 sky130_fd_sc_hd__a21oi_1 _1815_ (.A1(_0518_),
    .A2(_0695_),
    .B1(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__mux4_1 _1816_ (.A0(\RAM[72][1] ),
    .A1(\RAM[73][1] ),
    .A2(\RAM[74][1] ),
    .A3(\RAM[75][1] ),
    .S0(_0622_),
    .S1(_0618_),
    .X(_0699_));
 sky130_fd_sc_hd__o21ai_1 _1817_ (.A1(_0536_),
    .A2(_0699_),
    .B1(_0624_),
    .Y(_0700_));
 sky130_fd_sc_hd__o32a_1 _1818_ (.A1(_0624_),
    .A2(_0692_),
    .A3(_0694_),
    .B1(_0698_),
    .B2(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__mux4_1 _1819_ (.A0(\RAM[84][1] ),
    .A1(\RAM[85][1] ),
    .A2(\RAM[86][1] ),
    .A3(\RAM[87][1] ),
    .S0(_0520_),
    .S1(_0618_),
    .X(_0702_));
 sky130_fd_sc_hd__mux4_1 _1820_ (.A0(\RAM[88][1] ),
    .A1(\RAM[89][1] ),
    .A2(\RAM[90][1] ),
    .A3(\RAM[91][1] ),
    .S0(_0520_),
    .S1(_0618_),
    .X(_0703_));
 sky130_fd_sc_hd__a22o_1 _1821_ (.A1(_0627_),
    .A2(_0702_),
    .B1(_0703_),
    .B2(_0578_),
    .X(_0704_));
 sky130_fd_sc_hd__mux4_1 _1822_ (.A0(\RAM[92][1] ),
    .A1(\RAM[93][1] ),
    .A2(\RAM[94][1] ),
    .A3(\RAM[95][1] ),
    .S0(_0520_),
    .S1(_0618_),
    .X(_0705_));
 sky130_fd_sc_hd__mux4_1 _1823_ (.A0(\RAM[80][1] ),
    .A1(\RAM[81][1] ),
    .A2(\RAM[82][1] ),
    .A3(\RAM[83][1] ),
    .S0(_0528_),
    .S1(_0558_),
    .X(_0706_));
 sky130_fd_sc_hd__a22o_1 _1824_ (.A1(_0587_),
    .A2(_0705_),
    .B1(_0706_),
    .B2(_0634_),
    .X(_0707_));
 sky130_fd_sc_hd__nor2_1 _1825_ (.A(_0704_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__mux4_1 _1826_ (.A0(\RAM[104][1] ),
    .A1(\RAM[105][1] ),
    .A2(\RAM[106][1] ),
    .A3(\RAM[107][1] ),
    .S0(_0519_),
    .S1(_0548_),
    .X(_0709_));
 sky130_fd_sc_hd__or2_1 _1827_ (.A(_0535_),
    .B(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__mux4_1 _1828_ (.A0(\RAM[108][1] ),
    .A1(\RAM[109][1] ),
    .A2(\RAM[110][1] ),
    .A3(\RAM[111][1] ),
    .S0(_0519_),
    .S1(_0548_),
    .X(_0711_));
 sky130_fd_sc_hd__or2_1 _1829_ (.A(_0614_),
    .B(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__mux4_1 _1830_ (.A0(\RAM[100][1] ),
    .A1(\RAM[101][1] ),
    .A2(\RAM[102][1] ),
    .A3(\RAM[103][1] ),
    .S0(_0519_),
    .S1(_0548_),
    .X(_0713_));
 sky130_fd_sc_hd__mux4_1 _1831_ (.A0(\RAM[96][1] ),
    .A1(\RAM[97][1] ),
    .A2(\RAM[98][1] ),
    .A3(\RAM[99][1] ),
    .S0(_0519_),
    .S1(_0548_),
    .X(_0714_));
 sky130_fd_sc_hd__a22o_1 _1832_ (.A1(_0590_),
    .A2(_0713_),
    .B1(_0714_),
    .B2(_0584_),
    .X(_0715_));
 sky130_fd_sc_hd__a31o_1 _1833_ (.A1(_0624_),
    .A2(_0710_),
    .A3(_0712_),
    .B1(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__mux4_1 _1834_ (.A0(\RAM[112][1] ),
    .A1(\RAM[113][1] ),
    .A2(\RAM[114][1] ),
    .A3(\RAM[115][1] ),
    .S0(_0528_),
    .S1(_0558_),
    .X(_0717_));
 sky130_fd_sc_hd__mux4_1 _1835_ (.A0(\RAM[120][1] ),
    .A1(\RAM[121][1] ),
    .A2(\RAM[122][1] ),
    .A3(\RAM[123][1] ),
    .S0(_0527_),
    .S1(_0548_),
    .X(_0718_));
 sky130_fd_sc_hd__mux4_1 _1836_ (.A0(\RAM[124][1] ),
    .A1(\RAM[125][1] ),
    .A2(\RAM[126][1] ),
    .A3(\RAM[127][1] ),
    .S0(_0527_),
    .S1(_0566_),
    .X(_0719_));
 sky130_fd_sc_hd__o22a_1 _1837_ (.A1(_0561_),
    .A2(_0718_),
    .B1(_0719_),
    .B2(_0564_),
    .X(_0720_));
 sky130_fd_sc_hd__mux4_1 _1838_ (.A0(\RAM[116][1] ),
    .A1(\RAM[117][1] ),
    .A2(\RAM[118][1] ),
    .A3(\RAM[119][1] ),
    .S0(_0571_),
    .S1(_0595_),
    .X(_0721_));
 sky130_fd_sc_hd__o21ba_1 _1839_ (.A1(_0570_),
    .A2(_0721_),
    .B1_N(_0574_),
    .X(_0722_));
 sky130_fd_sc_hd__o211a_1 _1840_ (.A1(_0557_),
    .A2(_0717_),
    .B1(_0720_),
    .C1(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__a21oi_1 _1841_ (.A1(_0592_),
    .A2(_0716_),
    .B1(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__o221a_1 _1842_ (.A1(_0513_),
    .A2(_0701_),
    .B1(_0708_),
    .B2(_0602_),
    .C1(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__a22oi_4 _1843_ (.A1(_0667_),
    .A2(_0688_),
    .B1(_0725_),
    .B2(net7),
    .Y(net14));
 sky130_fd_sc_hd__mux4_1 _1844_ (.A0(\RAM[72][2] ),
    .A1(\RAM[73][2] ),
    .A2(\RAM[74][2] ),
    .A3(\RAM[75][2] ),
    .S0(_0637_),
    .S1(_0638_),
    .X(_0726_));
 sky130_fd_sc_hd__or2_1 _1845_ (.A(_0535_),
    .B(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _1846_ (.A0(\RAM[78][2] ),
    .A1(\RAM[79][2] ),
    .S(_0528_),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _1847_ (.A0(\RAM[76][2] ),
    .A1(\RAM[77][2] ),
    .S(_0565_),
    .X(_0729_));
 sky130_fd_sc_hd__a21o_1 _1848_ (.A1(_0524_),
    .A2(_0729_),
    .B1(_0614_),
    .X(_0730_));
 sky130_fd_sc_hd__a21o_1 _1849_ (.A1(_0550_),
    .A2(_0728_),
    .B1(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _1850_ (.A0(\RAM[68][2] ),
    .A1(\RAM[69][2] ),
    .S(_0528_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _1851_ (.A0(\RAM[70][2] ),
    .A1(\RAM[71][2] ),
    .S(_0519_),
    .X(_0733_));
 sky130_fd_sc_hd__and2_1 _1852_ (.A(_0549_),
    .B(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__a211o_1 _1853_ (.A1(_0525_),
    .A2(_0732_),
    .B1(_0734_),
    .C1(_0531_),
    .X(_0735_));
 sky130_fd_sc_hd__mux4_1 _1854_ (.A0(\RAM[64][2] ),
    .A1(\RAM[65][2] ),
    .A2(\RAM[66][2] ),
    .A3(\RAM[67][2] ),
    .S0(_0538_),
    .S1(_0628_),
    .X(_0736_));
 sky130_fd_sc_hd__o21ba_1 _1855_ (.A1(_0535_),
    .A2(_0736_),
    .B1_N(_0624_),
    .X(_0737_));
 sky130_fd_sc_hd__a32o_1 _1856_ (.A1(_0515_),
    .A2(_0727_),
    .A3(_0731_),
    .B1(_0735_),
    .B2(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__mux4_1 _1857_ (.A0(\RAM[84][2] ),
    .A1(\RAM[85][2] ),
    .A2(\RAM[86][2] ),
    .A3(\RAM[87][2] ),
    .S0(_0538_),
    .S1(_0628_),
    .X(_0739_));
 sky130_fd_sc_hd__mux4_1 _1858_ (.A0(\RAM[88][2] ),
    .A1(\RAM[89][2] ),
    .A2(\RAM[90][2] ),
    .A3(\RAM[91][2] ),
    .S0(_0622_),
    .S1(_0549_),
    .X(_0740_));
 sky130_fd_sc_hd__a22o_1 _1859_ (.A1(_0627_),
    .A2(_0739_),
    .B1(_0740_),
    .B2(_0578_),
    .X(_0741_));
 sky130_fd_sc_hd__mux4_1 _1860_ (.A0(\RAM[92][2] ),
    .A1(\RAM[93][2] ),
    .A2(\RAM[94][2] ),
    .A3(\RAM[95][2] ),
    .S0(_0538_),
    .S1(_0628_),
    .X(_0742_));
 sky130_fd_sc_hd__mux4_1 _1861_ (.A0(\RAM[80][2] ),
    .A1(\RAM[81][2] ),
    .A2(\RAM[82][2] ),
    .A3(\RAM[83][2] ),
    .S0(_0622_),
    .S1(_0549_),
    .X(_0743_));
 sky130_fd_sc_hd__a22o_1 _1862_ (.A1(_0587_),
    .A2(_0742_),
    .B1(_0743_),
    .B2(_0634_),
    .X(_0744_));
 sky130_fd_sc_hd__o21ba_1 _1863_ (.A1(_0741_),
    .A2(_0744_),
    .B1_N(_0602_),
    .X(_0745_));
 sky130_fd_sc_hd__mux4_1 _1864_ (.A0(\RAM[108][2] ),
    .A1(\RAM[109][2] ),
    .A2(\RAM[110][2] ),
    .A3(\RAM[111][2] ),
    .S0(_0543_),
    .S1(_0595_),
    .X(_0746_));
 sky130_fd_sc_hd__mux4_1 _1865_ (.A0(\RAM[104][2] ),
    .A1(\RAM[105][2] ),
    .A2(\RAM[106][2] ),
    .A3(\RAM[107][2] ),
    .S0(_0526_),
    .S1(net2),
    .X(_0747_));
 sky130_fd_sc_hd__or2_1 _1866_ (.A(_0534_),
    .B(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__o211a_1 _1867_ (.A1(_0614_),
    .A2(_0746_),
    .B1(_0748_),
    .C1(_0514_),
    .X(_0749_));
 sky130_fd_sc_hd__mux4_1 _1868_ (.A0(\RAM[96][2] ),
    .A1(\RAM[97][2] ),
    .A2(\RAM[98][2] ),
    .A3(\RAM[99][2] ),
    .S0(_0606_),
    .S1(_0608_),
    .X(_0750_));
 sky130_fd_sc_hd__mux4_1 _1869_ (.A0(\RAM[100][2] ),
    .A1(\RAM[101][2] ),
    .A2(\RAM[102][2] ),
    .A3(\RAM[103][2] ),
    .S0(_0606_),
    .S1(_0608_),
    .X(_0751_));
 sky130_fd_sc_hd__a22o_1 _1870_ (.A1(_0634_),
    .A2(_0750_),
    .B1(_0751_),
    .B2(_0627_),
    .X(_0752_));
 sky130_fd_sc_hd__mux4_1 _1871_ (.A0(\RAM[116][2] ),
    .A1(\RAM[117][2] ),
    .A2(\RAM[118][2] ),
    .A3(\RAM[119][2] ),
    .S0(_0537_),
    .S1(_0607_),
    .X(_0753_));
 sky130_fd_sc_hd__mux4_1 _1872_ (.A0(\RAM[120][2] ),
    .A1(\RAM[121][2] ),
    .A2(\RAM[122][2] ),
    .A3(\RAM[123][2] ),
    .S0(_0519_),
    .S1(_0607_),
    .X(_0754_));
 sky130_fd_sc_hd__o22a_1 _1873_ (.A1(_0569_),
    .A2(_0753_),
    .B1(_0754_),
    .B2(_0560_),
    .X(_0755_));
 sky130_fd_sc_hd__mux4_1 _1874_ (.A0(\RAM[124][2] ),
    .A1(\RAM[125][2] ),
    .A2(\RAM[126][2] ),
    .A3(\RAM[127][2] ),
    .S0(_0537_),
    .S1(_0607_),
    .X(_0756_));
 sky130_fd_sc_hd__mux4_1 _1875_ (.A0(\RAM[112][2] ),
    .A1(\RAM[113][2] ),
    .A2(\RAM[114][2] ),
    .A3(\RAM[115][2] ),
    .S0(_0537_),
    .S1(_0607_),
    .X(_0757_));
 sky130_fd_sc_hd__o22a_1 _1876_ (.A1(_0564_),
    .A2(_0756_),
    .B1(_0757_),
    .B2(_0556_),
    .X(_0758_));
 sky130_fd_sc_hd__a21bo_1 _1877_ (.A1(_0755_),
    .A2(_0758_),
    .B1_N(_0573_),
    .X(_0759_));
 sky130_fd_sc_hd__o311a_1 _1878_ (.A1(_0573_),
    .A2(_0749_),
    .A3(_0752_),
    .B1(_0759_),
    .C1(net6),
    .X(_0760_));
 sky130_fd_sc_hd__a211o_1 _1879_ (.A1(_0605_),
    .A2(_0738_),
    .B1(_0745_),
    .C1(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _1880_ (.A0(\RAM[6][2] ),
    .A1(\RAM[7][2] ),
    .S(_0521_),
    .X(_0762_));
 sky130_fd_sc_hd__mux2_1 _1881_ (.A0(\RAM[4][2] ),
    .A1(\RAM[5][2] ),
    .S(_0528_),
    .X(_0763_));
 sky130_fd_sc_hd__a21o_1 _1882_ (.A1(_0525_),
    .A2(_0763_),
    .B1(_0531_),
    .X(_0764_));
 sky130_fd_sc_hd__a21oi_1 _1883_ (.A1(_0518_),
    .A2(_0762_),
    .B1(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__mux4_1 _1884_ (.A0(\RAM[0][2] ),
    .A1(\RAM[1][2] ),
    .A2(\RAM[2][2] ),
    .A3(\RAM[3][2] ),
    .S0(_0539_),
    .S1(_0550_),
    .X(_0766_));
 sky130_fd_sc_hd__nor2_1 _1885_ (.A(_0536_),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__mux2_1 _1886_ (.A0(\RAM[14][2] ),
    .A1(\RAM[15][2] ),
    .S(_0521_),
    .X(_0768_));
 sky130_fd_sc_hd__mux2_1 _1887_ (.A0(\RAM[12][2] ),
    .A1(\RAM[13][2] ),
    .S(_0544_),
    .X(_0769_));
 sky130_fd_sc_hd__a21o_1 _1888_ (.A1(_0525_),
    .A2(_0769_),
    .B1(_0531_),
    .X(_0770_));
 sky130_fd_sc_hd__a21oi_1 _1889_ (.A1(_0518_),
    .A2(_0768_),
    .B1(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__mux4_1 _1890_ (.A0(\RAM[8][2] ),
    .A1(\RAM[9][2] ),
    .A2(\RAM[10][2] ),
    .A3(\RAM[11][2] ),
    .S0(_0539_),
    .S1(_0550_),
    .X(_0772_));
 sky130_fd_sc_hd__o21ai_1 _1891_ (.A1(_0536_),
    .A2(_0772_),
    .B1(_0515_),
    .Y(_0773_));
 sky130_fd_sc_hd__o32a_1 _1892_ (.A1(_0515_),
    .A2(_0765_),
    .A3(_0767_),
    .B1(_0771_),
    .B2(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__nor2_1 _1893_ (.A(_0513_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__mux4_1 _1894_ (.A0(\RAM[48][2] ),
    .A1(\RAM[49][2] ),
    .A2(\RAM[50][2] ),
    .A3(\RAM[51][2] ),
    .S0(_0611_),
    .S1(_0558_),
    .X(_0776_));
 sky130_fd_sc_hd__mux4_1 _1895_ (.A0(\RAM[56][2] ),
    .A1(\RAM[57][2] ),
    .A2(\RAM[58][2] ),
    .A3(\RAM[59][2] ),
    .S0(_0527_),
    .S1(_0566_),
    .X(_0777_));
 sky130_fd_sc_hd__mux4_1 _1896_ (.A0(\RAM[60][2] ),
    .A1(\RAM[61][2] ),
    .A2(\RAM[62][2] ),
    .A3(\RAM[63][2] ),
    .S0(_0565_),
    .S1(_0566_),
    .X(_0778_));
 sky130_fd_sc_hd__o22a_1 _1897_ (.A1(_0561_),
    .A2(_0777_),
    .B1(_0778_),
    .B2(_0564_),
    .X(_0779_));
 sky130_fd_sc_hd__mux4_1 _1898_ (.A0(\RAM[52][2] ),
    .A1(\RAM[53][2] ),
    .A2(\RAM[54][2] ),
    .A3(\RAM[55][2] ),
    .S0(_0543_),
    .S1(_0638_),
    .X(_0780_));
 sky130_fd_sc_hd__o21ba_1 _1899_ (.A1(_0570_),
    .A2(_0780_),
    .B1_N(_0574_),
    .X(_0781_));
 sky130_fd_sc_hd__o211a_1 _1900_ (.A1(_0557_),
    .A2(_0776_),
    .B1(_0779_),
    .C1(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__mux4_1 _1901_ (.A0(\RAM[36][2] ),
    .A1(\RAM[37][2] ),
    .A2(\RAM[38][2] ),
    .A3(\RAM[39][2] ),
    .S0(_0527_),
    .S1(_0566_),
    .X(_0783_));
 sky130_fd_sc_hd__mux4_1 _1902_ (.A0(\RAM[32][2] ),
    .A1(\RAM[33][2] ),
    .A2(\RAM[34][2] ),
    .A3(\RAM[35][2] ),
    .S0(_0543_),
    .S1(_0595_),
    .X(_0784_));
 sky130_fd_sc_hd__a22o_1 _1903_ (.A1(_0590_),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_0584_),
    .X(_0785_));
 sky130_fd_sc_hd__mux4_1 _1904_ (.A0(\RAM[44][2] ),
    .A1(\RAM[45][2] ),
    .A2(\RAM[46][2] ),
    .A3(\RAM[47][2] ),
    .S0(_0527_),
    .S1(_0566_),
    .X(_0786_));
 sky130_fd_sc_hd__mux4_1 _1905_ (.A0(\RAM[40][2] ),
    .A1(\RAM[41][2] ),
    .A2(\RAM[42][2] ),
    .A3(\RAM[43][2] ),
    .S0(_0526_),
    .S1(net2),
    .X(_0787_));
 sky130_fd_sc_hd__or2_1 _1906_ (.A(_0534_),
    .B(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__o211a_1 _1907_ (.A1(_0614_),
    .A2(_0786_),
    .B1(_0788_),
    .C1(_0514_),
    .X(_0789_));
 sky130_fd_sc_hd__o21a_1 _1908_ (.A1(_0785_),
    .A2(_0789_),
    .B1(_0592_),
    .X(_0790_));
 sky130_fd_sc_hd__mux4_1 _1909_ (.A0(\RAM[20][2] ),
    .A1(\RAM[21][2] ),
    .A2(\RAM[22][2] ),
    .A3(\RAM[23][2] ),
    .S0(_0571_),
    .S1(_0516_),
    .X(_0791_));
 sky130_fd_sc_hd__mux4_1 _1910_ (.A0(\RAM[24][2] ),
    .A1(\RAM[25][2] ),
    .A2(\RAM[26][2] ),
    .A3(\RAM[27][2] ),
    .S0(_0637_),
    .S1(_0638_),
    .X(_0792_));
 sky130_fd_sc_hd__a22o_1 _1911_ (.A1(_0627_),
    .A2(_0791_),
    .B1(_0792_),
    .B2(_0578_),
    .X(_0793_));
 sky130_fd_sc_hd__mux4_1 _1912_ (.A0(\RAM[28][2] ),
    .A1(\RAM[29][2] ),
    .A2(\RAM[30][2] ),
    .A3(\RAM[31][2] ),
    .S0(_0571_),
    .S1(_0595_),
    .X(_0794_));
 sky130_fd_sc_hd__mux4_1 _1913_ (.A0(\RAM[16][2] ),
    .A1(\RAM[17][2] ),
    .A2(\RAM[18][2] ),
    .A3(\RAM[19][2] ),
    .S0(_0637_),
    .S1(_0638_),
    .X(_0795_));
 sky130_fd_sc_hd__a22o_1 _1914_ (.A1(_0587_),
    .A2(_0794_),
    .B1(_0795_),
    .B2(_0634_),
    .X(_0796_));
 sky130_fd_sc_hd__o21ba_1 _1915_ (.A1(_0793_),
    .A2(_0796_),
    .B1_N(_0602_),
    .X(_0797_));
 sky130_fd_sc_hd__or4_1 _1916_ (.A(net7),
    .B(_0782_),
    .C(_0790_),
    .D(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__o22a_1 _1917_ (.A1(_0555_),
    .A2(_0761_),
    .B1(_0775_),
    .B2(_0798_),
    .X(net15));
 sky130_fd_sc_hd__mux2_1 _1918_ (.A0(\RAM[70][3] ),
    .A1(\RAM[71][3] ),
    .S(_0544_),
    .X(_0799_));
 sky130_fd_sc_hd__mux2_1 _1919_ (.A0(\RAM[68][3] ),
    .A1(\RAM[69][3] ),
    .S(_0606_),
    .X(_0800_));
 sky130_fd_sc_hd__a21o_1 _1920_ (.A1(_0524_),
    .A2(_0800_),
    .B1(_0614_),
    .X(_0801_));
 sky130_fd_sc_hd__a21oi_1 _1921_ (.A1(_0518_),
    .A2(_0799_),
    .B1(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__mux4_1 _1922_ (.A0(\RAM[64][3] ),
    .A1(\RAM[65][3] ),
    .A2(\RAM[66][3] ),
    .A3(\RAM[67][3] ),
    .S0(_0528_),
    .S1(_0558_),
    .X(_0803_));
 sky130_fd_sc_hd__nor2_1 _1923_ (.A(_0536_),
    .B(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__mux2_1 _1924_ (.A0(\RAM[78][3] ),
    .A1(\RAM[79][3] ),
    .S(_0539_),
    .X(_0805_));
 sky130_fd_sc_hd__mux2_1 _1925_ (.A0(\RAM[76][3] ),
    .A1(\RAM[77][3] ),
    .S(_0622_),
    .X(_0806_));
 sky130_fd_sc_hd__a21o_1 _1926_ (.A1(_0525_),
    .A2(_0806_),
    .B1(_0531_),
    .X(_0807_));
 sky130_fd_sc_hd__a21oi_1 _1927_ (.A1(_0518_),
    .A2(_0805_),
    .B1(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__mux4_1 _1928_ (.A0(\RAM[72][3] ),
    .A1(\RAM[73][3] ),
    .A2(\RAM[74][3] ),
    .A3(\RAM[75][3] ),
    .S0(_0611_),
    .S1(_0517_),
    .X(_0809_));
 sky130_fd_sc_hd__o21ai_1 _1929_ (.A1(_0536_),
    .A2(_0809_),
    .B1(_0515_),
    .Y(_0810_));
 sky130_fd_sc_hd__o32a_1 _1930_ (.A1(_0515_),
    .A2(_0802_),
    .A3(_0804_),
    .B1(_0808_),
    .B2(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__mux4_1 _1931_ (.A0(\RAM[84][3] ),
    .A1(\RAM[85][3] ),
    .A2(\RAM[86][3] ),
    .A3(\RAM[87][3] ),
    .S0(_0611_),
    .S1(_0517_),
    .X(_0812_));
 sky130_fd_sc_hd__mux4_1 _1932_ (.A0(\RAM[88][3] ),
    .A1(\RAM[89][3] ),
    .A2(\RAM[90][3] ),
    .A3(\RAM[91][3] ),
    .S0(_0544_),
    .S1(_0517_),
    .X(_0813_));
 sky130_fd_sc_hd__a22o_1 _1933_ (.A1(_0627_),
    .A2(_0812_),
    .B1(_0813_),
    .B2(_0578_),
    .X(_0814_));
 sky130_fd_sc_hd__mux4_1 _1934_ (.A0(\RAM[92][3] ),
    .A1(\RAM[93][3] ),
    .A2(\RAM[94][3] ),
    .A3(\RAM[95][3] ),
    .S0(_0544_),
    .S1(_0517_),
    .X(_0815_));
 sky130_fd_sc_hd__mux4_1 _1935_ (.A0(\RAM[80][3] ),
    .A1(\RAM[81][3] ),
    .A2(\RAM[82][3] ),
    .A3(\RAM[83][3] ),
    .S0(_0544_),
    .S1(_0517_),
    .X(_0816_));
 sky130_fd_sc_hd__a22o_1 _1936_ (.A1(_0587_),
    .A2(_0815_),
    .B1(_0816_),
    .B2(_0634_),
    .X(_0817_));
 sky130_fd_sc_hd__nor2_1 _1937_ (.A(_0814_),
    .B(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__mux4_1 _1938_ (.A0(\RAM[104][3] ),
    .A1(\RAM[105][3] ),
    .A2(\RAM[106][3] ),
    .A3(\RAM[107][3] ),
    .S0(_0606_),
    .S1(_0608_),
    .X(_0819_));
 sky130_fd_sc_hd__o21a_1 _1939_ (.A1(_0535_),
    .A2(_0819_),
    .B1(_0624_),
    .X(_0820_));
 sky130_fd_sc_hd__mux4_1 _1940_ (.A0(\RAM[108][3] ),
    .A1(\RAM[109][3] ),
    .A2(\RAM[110][3] ),
    .A3(\RAM[111][3] ),
    .S0(_0571_),
    .S1(_0516_),
    .X(_0821_));
 sky130_fd_sc_hd__or2_1 _1941_ (.A(_0614_),
    .B(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__mux4_1 _1942_ (.A0(\RAM[100][3] ),
    .A1(\RAM[101][3] ),
    .A2(\RAM[102][3] ),
    .A3(\RAM[103][3] ),
    .S0(_0543_),
    .S1(_0595_),
    .X(_0823_));
 sky130_fd_sc_hd__mux4_1 _1943_ (.A0(\RAM[96][3] ),
    .A1(\RAM[97][3] ),
    .A2(\RAM[98][3] ),
    .A3(\RAM[99][3] ),
    .S0(_0606_),
    .S1(_0608_),
    .X(_0824_));
 sky130_fd_sc_hd__a22o_1 _1944_ (.A1(_0627_),
    .A2(_0823_),
    .B1(_0824_),
    .B2(_0634_),
    .X(_0825_));
 sky130_fd_sc_hd__a21o_1 _1945_ (.A1(_0820_),
    .A2(_0822_),
    .B1(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__mux4_1 _1946_ (.A0(\RAM[112][3] ),
    .A1(\RAM[113][3] ),
    .A2(\RAM[114][3] ),
    .A3(\RAM[115][3] ),
    .S0(_0544_),
    .S1(_0517_),
    .X(_0827_));
 sky130_fd_sc_hd__mux4_1 _1947_ (.A0(\RAM[120][3] ),
    .A1(\RAM[121][3] ),
    .A2(\RAM[122][3] ),
    .A3(\RAM[123][3] ),
    .S0(_0637_),
    .S1(_0638_),
    .X(_0828_));
 sky130_fd_sc_hd__mux4_1 _1948_ (.A0(\RAM[124][3] ),
    .A1(\RAM[125][3] ),
    .A2(\RAM[126][3] ),
    .A3(\RAM[127][3] ),
    .S0(_0637_),
    .S1(_0608_),
    .X(_0829_));
 sky130_fd_sc_hd__o22a_1 _1949_ (.A1(_0561_),
    .A2(_0828_),
    .B1(_0829_),
    .B2(_0564_),
    .X(_0830_));
 sky130_fd_sc_hd__mux4_1 _1950_ (.A0(\RAM[116][3] ),
    .A1(\RAM[117][3] ),
    .A2(\RAM[118][3] ),
    .A3(\RAM[119][3] ),
    .S0(_0538_),
    .S1(_0628_),
    .X(_0831_));
 sky130_fd_sc_hd__o21ba_1 _1951_ (.A1(_0570_),
    .A2(_0831_),
    .B1_N(_0574_),
    .X(_0832_));
 sky130_fd_sc_hd__o211a_1 _1952_ (.A1(_0557_),
    .A2(_0827_),
    .B1(_0830_),
    .C1(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__a21oi_1 _1953_ (.A1(_0592_),
    .A2(_0826_),
    .B1(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__o221a_1 _1954_ (.A1(_0513_),
    .A2(_0811_),
    .B1(_0818_),
    .B2(_0602_),
    .C1(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _1955_ (.A0(\RAM[6][3] ),
    .A1(\RAM[7][3] ),
    .S(_0521_),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_1 _1956_ (.A0(\RAM[4][3] ),
    .A1(\RAM[5][3] ),
    .S(_0611_),
    .X(_0837_));
 sky130_fd_sc_hd__a21o_1 _1957_ (.A1(_0525_),
    .A2(_0837_),
    .B1(_0531_),
    .X(_0838_));
 sky130_fd_sc_hd__a21oi_1 _1958_ (.A1(_0518_),
    .A2(_0836_),
    .B1(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__mux4_1 _1959_ (.A0(\RAM[0][3] ),
    .A1(\RAM[1][3] ),
    .A2(\RAM[2][3] ),
    .A3(\RAM[3][3] ),
    .S0(_0539_),
    .S1(_0550_),
    .X(_0840_));
 sky130_fd_sc_hd__nor2_1 _1960_ (.A(_0536_),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__mux2_1 _1961_ (.A0(\RAM[14][3] ),
    .A1(\RAM[15][3] ),
    .S(_0521_),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_1 _1962_ (.A0(\RAM[12][3] ),
    .A1(\RAM[13][3] ),
    .S(_0544_),
    .X(_0843_));
 sky130_fd_sc_hd__a21o_1 _1963_ (.A1(_0525_),
    .A2(_0843_),
    .B1(_0531_),
    .X(_0844_));
 sky130_fd_sc_hd__a21oi_1 _1964_ (.A1(_0518_),
    .A2(_0842_),
    .B1(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__mux4_1 _1965_ (.A0(\RAM[8][3] ),
    .A1(\RAM[9][3] ),
    .A2(\RAM[10][3] ),
    .A3(\RAM[11][3] ),
    .S0(_0521_),
    .S1(_0550_),
    .X(_0846_));
 sky130_fd_sc_hd__o21ai_1 _1966_ (.A1(_0536_),
    .A2(_0846_),
    .B1(_0515_),
    .Y(_0847_));
 sky130_fd_sc_hd__o32a_1 _1967_ (.A1(_0515_),
    .A2(_0839_),
    .A3(_0841_),
    .B1(_0845_),
    .B2(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__nor2_1 _1968_ (.A(_0513_),
    .B(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__mux4_1 _1969_ (.A0(\RAM[48][3] ),
    .A1(\RAM[49][3] ),
    .A2(\RAM[50][3] ),
    .A3(\RAM[51][3] ),
    .S0(_0611_),
    .S1(_0517_),
    .X(_0850_));
 sky130_fd_sc_hd__mux4_1 _1970_ (.A0(\RAM[56][3] ),
    .A1(\RAM[57][3] ),
    .A2(\RAM[58][3] ),
    .A3(\RAM[59][3] ),
    .S0(_0527_),
    .S1(_0566_),
    .X(_0851_));
 sky130_fd_sc_hd__mux4_1 _1971_ (.A0(\RAM[60][3] ),
    .A1(\RAM[61][3] ),
    .A2(\RAM[62][3] ),
    .A3(\RAM[63][3] ),
    .S0(_0571_),
    .S1(_0516_),
    .X(_0852_));
 sky130_fd_sc_hd__o22a_1 _1972_ (.A1(_0561_),
    .A2(_0851_),
    .B1(_0852_),
    .B2(_0564_),
    .X(_0853_));
 sky130_fd_sc_hd__mux4_1 _1973_ (.A0(\RAM[52][3] ),
    .A1(\RAM[53][3] ),
    .A2(\RAM[54][3] ),
    .A3(\RAM[55][3] ),
    .S0(_0637_),
    .S1(_0638_),
    .X(_0854_));
 sky130_fd_sc_hd__o21ba_1 _1974_ (.A1(_0570_),
    .A2(_0854_),
    .B1_N(_0574_),
    .X(_0855_));
 sky130_fd_sc_hd__o211a_1 _1975_ (.A1(_0557_),
    .A2(_0850_),
    .B1(_0853_),
    .C1(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__mux2_1 _1976_ (.A0(\RAM[40][3] ),
    .A1(\RAM[41][3] ),
    .S(_0537_),
    .X(_0857_));
 sky130_fd_sc_hd__or2_1 _1977_ (.A(_0638_),
    .B(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__mux2_1 _1978_ (.A0(\RAM[42][3] ),
    .A1(\RAM[43][3] ),
    .S(_0537_),
    .X(_0859_));
 sky130_fd_sc_hd__or2_1 _1979_ (.A(_0523_),
    .B(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__mux4_1 _1980_ (.A0(\RAM[32][3] ),
    .A1(\RAM[33][3] ),
    .A2(\RAM[34][3] ),
    .A3(\RAM[35][3] ),
    .S0(_0543_),
    .S1(_0595_),
    .X(_0861_));
 sky130_fd_sc_hd__a32o_1 _1981_ (.A1(_0578_),
    .A2(_0858_),
    .A3(_0860_),
    .B1(_0861_),
    .B2(_0584_),
    .X(_0862_));
 sky130_fd_sc_hd__mux4_1 _1982_ (.A0(\RAM[44][3] ),
    .A1(\RAM[45][3] ),
    .A2(\RAM[46][3] ),
    .A3(\RAM[47][3] ),
    .S0(_0571_),
    .S1(_0516_),
    .X(_0863_));
 sky130_fd_sc_hd__mux4_1 _1983_ (.A0(\RAM[36][3] ),
    .A1(\RAM[37][3] ),
    .A2(\RAM[38][3] ),
    .A3(\RAM[39][3] ),
    .S0(_0543_),
    .S1(_0638_),
    .X(_0864_));
 sky130_fd_sc_hd__a22o_1 _1984_ (.A1(_0587_),
    .A2(_0863_),
    .B1(_0864_),
    .B2(_0590_),
    .X(_0865_));
 sky130_fd_sc_hd__o21a_1 _1985_ (.A1(_0862_),
    .A2(_0865_),
    .B1(_0592_),
    .X(_0866_));
 sky130_fd_sc_hd__mux4_1 _1986_ (.A0(\RAM[20][3] ),
    .A1(\RAM[21][3] ),
    .A2(\RAM[22][3] ),
    .A3(\RAM[23][3] ),
    .S0(_0571_),
    .S1(_0595_),
    .X(_0867_));
 sky130_fd_sc_hd__mux4_1 _1987_ (.A0(\RAM[24][3] ),
    .A1(\RAM[25][3] ),
    .A2(\RAM[26][3] ),
    .A3(\RAM[27][3] ),
    .S0(_0637_),
    .S1(_0638_),
    .X(_0868_));
 sky130_fd_sc_hd__a22o_1 _1988_ (.A1(_0627_),
    .A2(_0867_),
    .B1(_0868_),
    .B2(_0578_),
    .X(_0869_));
 sky130_fd_sc_hd__mux4_1 _1989_ (.A0(\RAM[28][3] ),
    .A1(\RAM[29][3] ),
    .A2(\RAM[30][3] ),
    .A3(\RAM[31][3] ),
    .S0(_0543_),
    .S1(_0595_),
    .X(_0870_));
 sky130_fd_sc_hd__mux4_1 _1990_ (.A0(\RAM[16][3] ),
    .A1(\RAM[17][3] ),
    .A2(\RAM[18][3] ),
    .A3(\RAM[19][3] ),
    .S0(_0637_),
    .S1(_0608_),
    .X(_0871_));
 sky130_fd_sc_hd__a22o_1 _1991_ (.A1(_0587_),
    .A2(_0870_),
    .B1(_0871_),
    .B2(_0634_),
    .X(_0872_));
 sky130_fd_sc_hd__o21ba_1 _1992_ (.A1(_0869_),
    .A2(_0872_),
    .B1_N(_0602_),
    .X(_0873_));
 sky130_fd_sc_hd__or4_1 _1993_ (.A(net7),
    .B(_0856_),
    .C(_0866_),
    .D(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__o2bb2a_1 _1994_ (.A1_N(net7),
    .A2_N(_0835_),
    .B1(_0849_),
    .B2(_0874_),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 _1995_ (.A(net8),
    .X(_0875_));
 sky130_fd_sc_hd__clkbuf_4 _1996_ (.A(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__nand2_4 _1997_ (.A(_0520_),
    .B(_0523_),
    .Y(_0877_));
 sky130_fd_sc_hd__or2_4 _1998_ (.A(_0570_),
    .B(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__nand2_8 _1999_ (.A(net7),
    .B(net12),
    .Y(_0879_));
 sky130_fd_sc_hd__or2_1 _2000_ (.A(_0513_),
    .B(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__buf_4 _2001_ (.A(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__nor2_2 _2002_ (.A(_0878_),
    .B(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__mux2_1 _2003_ (.A0(\RAM[69][0] ),
    .A1(_0876_),
    .S(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__clkbuf_1 _2004_ (.A(_0883_),
    .X(_0000_));
 sky130_fd_sc_hd__clkbuf_4 _2005_ (.A(net9),
    .X(_0884_));
 sky130_fd_sc_hd__buf_4 _2006_ (.A(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _2007_ (.A0(\RAM[69][1] ),
    .A1(_0885_),
    .S(_0882_),
    .X(_0886_));
 sky130_fd_sc_hd__clkbuf_1 _2008_ (.A(_0886_),
    .X(_0001_));
 sky130_fd_sc_hd__clkbuf_4 _2009_ (.A(net10),
    .X(_0887_));
 sky130_fd_sc_hd__clkbuf_4 _2010_ (.A(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _2011_ (.A0(\RAM[69][2] ),
    .A1(_0888_),
    .S(_0882_),
    .X(_0889_));
 sky130_fd_sc_hd__clkbuf_1 _2012_ (.A(_0889_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_4 _2013_ (.A(net11),
    .X(_0890_));
 sky130_fd_sc_hd__buf_4 _2014_ (.A(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_1 _2015_ (.A0(\RAM[69][3] ),
    .A1(_0891_),
    .S(_0882_),
    .X(_0892_));
 sky130_fd_sc_hd__clkbuf_1 _2016_ (.A(_0892_),
    .X(_0003_));
 sky130_fd_sc_hd__buf_4 _2017_ (.A(_0875_),
    .X(_0893_));
 sky130_fd_sc_hd__nor2_4 _2018_ (.A(_0877_),
    .B(_0561_),
    .Y(_0894_));
 sky130_fd_sc_hd__nor2_4 _2019_ (.A(_0602_),
    .B(_0879_),
    .Y(_0895_));
 sky130_fd_sc_hd__nand2_2 _2020_ (.A(_0894_),
    .B(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__mux2_1 _2021_ (.A0(_0893_),
    .A1(\RAM[89][0] ),
    .S(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__clkbuf_1 _2022_ (.A(_0897_),
    .X(_0004_));
 sky130_fd_sc_hd__buf_6 _2023_ (.A(_0884_),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _2024_ (.A0(_0898_),
    .A1(\RAM[89][1] ),
    .S(_0896_),
    .X(_0899_));
 sky130_fd_sc_hd__clkbuf_1 _2025_ (.A(_0899_),
    .X(_0005_));
 sky130_fd_sc_hd__buf_4 _2026_ (.A(_0887_),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _2027_ (.A0(_0900_),
    .A1(\RAM[89][2] ),
    .S(_0896_),
    .X(_0901_));
 sky130_fd_sc_hd__clkbuf_1 _2028_ (.A(_0901_),
    .X(_0006_));
 sky130_fd_sc_hd__buf_4 _2029_ (.A(_0890_),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_1 _2030_ (.A0(_0902_),
    .A1(\RAM[89][3] ),
    .S(_0896_),
    .X(_0903_));
 sky130_fd_sc_hd__clkbuf_1 _2031_ (.A(_0903_),
    .X(_0007_));
 sky130_fd_sc_hd__nand2_8 _2032_ (.A(_0544_),
    .B(_0618_),
    .Y(_0904_));
 sky130_fd_sc_hd__nor2_8 _2033_ (.A(_0904_),
    .B(_0561_),
    .Y(_0905_));
 sky130_fd_sc_hd__nand2b_4 _2034_ (.A_N(net7),
    .B(net12),
    .Y(_0906_));
 sky130_fd_sc_hd__nor2_4 _2035_ (.A(_0574_),
    .B(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__nand2_1 _2036_ (.A(_0905_),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__mux2_1 _2037_ (.A0(_0893_),
    .A1(\RAM[59][0] ),
    .S(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__clkbuf_1 _2038_ (.A(_0909_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _2039_ (.A0(_0898_),
    .A1(\RAM[59][1] ),
    .S(_0908_),
    .X(_0910_));
 sky130_fd_sc_hd__clkbuf_1 _2040_ (.A(_0910_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _2041_ (.A0(_0900_),
    .A1(\RAM[59][2] ),
    .S(_0908_),
    .X(_0911_));
 sky130_fd_sc_hd__clkbuf_1 _2042_ (.A(_0911_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _2043_ (.A0(_0902_),
    .A1(\RAM[59][3] ),
    .S(_0908_),
    .X(_0912_));
 sky130_fd_sc_hd__clkbuf_1 _2044_ (.A(_0912_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _2045_ (.A(_0574_),
    .B(_0906_),
    .X(_0913_));
 sky130_fd_sc_hd__clkbuf_4 _2046_ (.A(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__or2_1 _2047_ (.A(_0877_),
    .B(_0557_),
    .X(_0915_));
 sky130_fd_sc_hd__buf_6 _2048_ (.A(_0915_),
    .X(_0916_));
 sky130_fd_sc_hd__nor2_2 _2049_ (.A(_0914_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__mux2_1 _2050_ (.A0(\RAM[49][0] ),
    .A1(_0876_),
    .S(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__clkbuf_1 _2051_ (.A(_0918_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _2052_ (.A0(\RAM[49][1] ),
    .A1(_0885_),
    .S(_0917_),
    .X(_0919_));
 sky130_fd_sc_hd__clkbuf_1 _2053_ (.A(_0919_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _2054_ (.A0(\RAM[49][2] ),
    .A1(_0888_),
    .S(_0917_),
    .X(_0920_));
 sky130_fd_sc_hd__clkbuf_1 _2055_ (.A(_0920_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _2056_ (.A0(\RAM[49][3] ),
    .A1(_0891_),
    .S(_0917_),
    .X(_0921_));
 sky130_fd_sc_hd__clkbuf_1 _2057_ (.A(_0921_),
    .X(_0015_));
 sky130_fd_sc_hd__nor2_8 _2058_ (.A(_0570_),
    .B(_0904_),
    .Y(_0922_));
 sky130_fd_sc_hd__or2b_2 _2059_ (.A(net5),
    .B_N(net6),
    .X(_0923_));
 sky130_fd_sc_hd__nor2_2 _2060_ (.A(_0923_),
    .B(_0906_),
    .Y(_0924_));
 sky130_fd_sc_hd__nand2_2 _2061_ (.A(_0922_),
    .B(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__mux2_1 _2062_ (.A0(_0893_),
    .A1(\RAM[39][0] ),
    .S(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__clkbuf_1 _2063_ (.A(_0926_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _2064_ (.A0(_0898_),
    .A1(\RAM[39][1] ),
    .S(_0925_),
    .X(_0927_));
 sky130_fd_sc_hd__clkbuf_1 _2065_ (.A(_0927_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _2066_ (.A0(_0900_),
    .A1(\RAM[39][2] ),
    .S(_0925_),
    .X(_0928_));
 sky130_fd_sc_hd__clkbuf_1 _2067_ (.A(_0928_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _2068_ (.A0(_0902_),
    .A1(\RAM[39][3] ),
    .S(_0925_),
    .X(_0929_));
 sky130_fd_sc_hd__clkbuf_1 _2069_ (.A(_0929_),
    .X(_0019_));
 sky130_fd_sc_hd__or2_4 _2070_ (.A(_0904_),
    .B(_0557_),
    .X(_0930_));
 sky130_fd_sc_hd__or2_1 _2071_ (.A(_0601_),
    .B(_0906_),
    .X(_0931_));
 sky130_fd_sc_hd__buf_4 _2072_ (.A(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__nor2_2 _2073_ (.A(_0930_),
    .B(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__mux2_1 _2074_ (.A0(\RAM[19][0] ),
    .A1(_0876_),
    .S(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__clkbuf_1 _2075_ (.A(_0934_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _2076_ (.A0(\RAM[19][1] ),
    .A1(_0885_),
    .S(_0933_),
    .X(_0935_));
 sky130_fd_sc_hd__clkbuf_1 _2077_ (.A(_0935_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _2078_ (.A0(\RAM[19][2] ),
    .A1(_0888_),
    .S(_0933_),
    .X(_0936_));
 sky130_fd_sc_hd__clkbuf_1 _2079_ (.A(_0936_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _2080_ (.A0(\RAM[19][3] ),
    .A1(_0891_),
    .S(_0933_),
    .X(_0937_));
 sky130_fd_sc_hd__clkbuf_1 _2081_ (.A(_0937_),
    .X(_0023_));
 sky130_fd_sc_hd__nor2_2 _2082_ (.A(_0513_),
    .B(_0879_),
    .Y(_0938_));
 sky130_fd_sc_hd__nor2_8 _2083_ (.A(_0904_),
    .B(_0564_),
    .Y(_0939_));
 sky130_fd_sc_hd__nand2_2 _2084_ (.A(_0938_),
    .B(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__mux2_1 _2085_ (.A0(_0893_),
    .A1(\RAM[79][0] ),
    .S(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__clkbuf_1 _2086_ (.A(_0941_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _2087_ (.A0(_0898_),
    .A1(\RAM[79][1] ),
    .S(_0940_),
    .X(_0942_));
 sky130_fd_sc_hd__clkbuf_1 _2088_ (.A(_0942_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _2089_ (.A0(_0900_),
    .A1(\RAM[79][2] ),
    .S(_0940_),
    .X(_0943_));
 sky130_fd_sc_hd__clkbuf_1 _2090_ (.A(_0943_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _2091_ (.A0(_0902_),
    .A1(\RAM[79][3] ),
    .S(_0940_),
    .X(_0944_));
 sky130_fd_sc_hd__clkbuf_1 _2092_ (.A(_0944_),
    .X(_0027_));
 sky130_fd_sc_hd__nor2_2 _2093_ (.A(_0602_),
    .B(_0906_),
    .Y(_0945_));
 sky130_fd_sc_hd__nor2_8 _2094_ (.A(_0877_),
    .B(_0564_),
    .Y(_0946_));
 sky130_fd_sc_hd__nand2_2 _2095_ (.A(_0945_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__mux2_1 _2096_ (.A0(_0893_),
    .A1(\RAM[29][0] ),
    .S(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__clkbuf_1 _2097_ (.A(_0948_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _2098_ (.A0(_0898_),
    .A1(\RAM[29][1] ),
    .S(_0947_),
    .X(_0949_));
 sky130_fd_sc_hd__clkbuf_1 _2099_ (.A(_0949_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _2100_ (.A0(_0900_),
    .A1(\RAM[29][2] ),
    .S(_0947_),
    .X(_0950_));
 sky130_fd_sc_hd__clkbuf_1 _2101_ (.A(_0950_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _2102_ (.A0(_0902_),
    .A1(\RAM[29][3] ),
    .S(_0947_),
    .X(_0951_));
 sky130_fd_sc_hd__clkbuf_1 _2103_ (.A(_0951_),
    .X(_0031_));
 sky130_fd_sc_hd__nor2_4 _2104_ (.A(_0904_),
    .B(_0557_),
    .Y(_0952_));
 sky130_fd_sc_hd__nor2_4 _2105_ (.A(_0923_),
    .B(_0879_),
    .Y(_0953_));
 sky130_fd_sc_hd__nand2_2 _2106_ (.A(_0952_),
    .B(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__mux2_1 _2107_ (.A0(_0893_),
    .A1(\RAM[99][0] ),
    .S(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__clkbuf_1 _2108_ (.A(_0955_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2109_ (.A0(_0898_),
    .A1(\RAM[99][1] ),
    .S(_0954_),
    .X(_0956_));
 sky130_fd_sc_hd__clkbuf_1 _2110_ (.A(_0956_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _2111_ (.A0(_0900_),
    .A1(\RAM[99][2] ),
    .S(_0954_),
    .X(_0957_));
 sky130_fd_sc_hd__clkbuf_1 _2112_ (.A(_0957_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2113_ (.A0(_0902_),
    .A1(\RAM[99][3] ),
    .S(_0954_),
    .X(_0958_));
 sky130_fd_sc_hd__clkbuf_1 _2114_ (.A(_0958_),
    .X(_0035_));
 sky130_fd_sc_hd__nand2_2 _2115_ (.A(_0946_),
    .B(_0953_),
    .Y(_0959_));
 sky130_fd_sc_hd__mux2_1 _2116_ (.A0(_0893_),
    .A1(\RAM[109][0] ),
    .S(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__clkbuf_1 _2117_ (.A(_0960_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2118_ (.A0(_0898_),
    .A1(\RAM[109][1] ),
    .S(_0959_),
    .X(_0961_));
 sky130_fd_sc_hd__clkbuf_1 _2119_ (.A(_0961_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2120_ (.A0(_0900_),
    .A1(\RAM[109][2] ),
    .S(_0959_),
    .X(_0962_));
 sky130_fd_sc_hd__clkbuf_1 _2121_ (.A(_0962_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2122_ (.A0(_0902_),
    .A1(\RAM[109][3] ),
    .S(_0959_),
    .X(_0963_));
 sky130_fd_sc_hd__clkbuf_1 _2123_ (.A(_0963_),
    .X(_0039_));
 sky130_fd_sc_hd__nor2_4 _2124_ (.A(_0574_),
    .B(_0879_),
    .Y(_0964_));
 sky130_fd_sc_hd__nand2_2 _2125_ (.A(_0922_),
    .B(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__mux2_1 _2126_ (.A0(_0893_),
    .A1(\RAM[119][0] ),
    .S(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__clkbuf_1 _2127_ (.A(_0966_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2128_ (.A0(_0898_),
    .A1(\RAM[119][1] ),
    .S(_0965_),
    .X(_0967_));
 sky130_fd_sc_hd__clkbuf_1 _2129_ (.A(_0967_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _2130_ (.A0(_0900_),
    .A1(\RAM[119][2] ),
    .S(_0965_),
    .X(_0968_));
 sky130_fd_sc_hd__clkbuf_1 _2131_ (.A(_0968_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _2132_ (.A0(_0902_),
    .A1(\RAM[119][3] ),
    .S(_0965_),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_1 _2133_ (.A(_0969_),
    .X(_0043_));
 sky130_fd_sc_hd__nand2_2 _2134_ (.A(_0939_),
    .B(_0964_),
    .Y(_0970_));
 sky130_fd_sc_hd__mux2_1 _2135_ (.A0(_0893_),
    .A1(\RAM[127][0] ),
    .S(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__clkbuf_1 _2136_ (.A(_0971_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _2137_ (.A0(_0898_),
    .A1(\RAM[127][1] ),
    .S(_0970_),
    .X(_0972_));
 sky130_fd_sc_hd__clkbuf_1 _2138_ (.A(_0972_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2139_ (.A0(_0900_),
    .A1(\RAM[127][2] ),
    .S(_0970_),
    .X(_0973_));
 sky130_fd_sc_hd__clkbuf_1 _2140_ (.A(_0973_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2141_ (.A0(_0902_),
    .A1(\RAM[127][3] ),
    .S(_0970_),
    .X(_0974_));
 sky130_fd_sc_hd__clkbuf_1 _2142_ (.A(_0974_),
    .X(_0047_));
 sky130_fd_sc_hd__or3_1 _2143_ (.A(_0611_),
    .B(_0608_),
    .C(_0563_),
    .X(_0975_));
 sky130_fd_sc_hd__buf_4 _2144_ (.A(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__or2_1 _2145_ (.A(_0513_),
    .B(_0906_),
    .X(_0977_));
 sky130_fd_sc_hd__buf_4 _2146_ (.A(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__nor2_2 _2147_ (.A(_0976_),
    .B(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__mux2_1 _2148_ (.A0(\RAM[12][0] ),
    .A1(_0876_),
    .S(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_1 _2149_ (.A(_0980_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _2150_ (.A0(\RAM[12][1] ),
    .A1(_0885_),
    .S(_0979_),
    .X(_0981_));
 sky130_fd_sc_hd__clkbuf_1 _2151_ (.A(_0981_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _2152_ (.A0(\RAM[12][2] ),
    .A1(_0888_),
    .S(_0979_),
    .X(_0982_));
 sky130_fd_sc_hd__clkbuf_1 _2153_ (.A(_0982_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _2154_ (.A0(\RAM[12][3] ),
    .A1(_0891_),
    .S(_0979_),
    .X(_0983_));
 sky130_fd_sc_hd__clkbuf_1 _2155_ (.A(_0983_),
    .X(_0051_));
 sky130_fd_sc_hd__nor2_2 _2156_ (.A(_0513_),
    .B(_0906_),
    .Y(_0984_));
 sky130_fd_sc_hd__nand2_2 _2157_ (.A(_0946_),
    .B(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__mux2_1 _2158_ (.A0(_0893_),
    .A1(\RAM[13][0] ),
    .S(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__clkbuf_1 _2159_ (.A(_0986_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _2160_ (.A0(_0898_),
    .A1(\RAM[13][1] ),
    .S(_0985_),
    .X(_0987_));
 sky130_fd_sc_hd__clkbuf_1 _2161_ (.A(_0987_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _2162_ (.A0(_0900_),
    .A1(\RAM[13][2] ),
    .S(_0985_),
    .X(_0988_));
 sky130_fd_sc_hd__clkbuf_1 _2163_ (.A(_0988_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2164_ (.A0(_0902_),
    .A1(\RAM[13][3] ),
    .S(_0985_),
    .X(_0989_));
 sky130_fd_sc_hd__clkbuf_1 _2165_ (.A(_0989_),
    .X(_0055_));
 sky130_fd_sc_hd__buf_4 _2166_ (.A(_0875_),
    .X(_0990_));
 sky130_fd_sc_hd__and3b_1 _2167_ (.A_N(_0521_),
    .B(_0517_),
    .C(_0586_),
    .X(_0991_));
 sky130_fd_sc_hd__buf_6 _2168_ (.A(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__nand2_2 _2169_ (.A(_0984_),
    .B(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__mux2_1 _2170_ (.A0(_0990_),
    .A1(\RAM[14][0] ),
    .S(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__clkbuf_1 _2171_ (.A(_0994_),
    .X(_0056_));
 sky130_fd_sc_hd__buf_4 _2172_ (.A(_0884_),
    .X(_0995_));
 sky130_fd_sc_hd__mux2_1 _2173_ (.A0(_0995_),
    .A1(\RAM[14][1] ),
    .S(_0993_),
    .X(_0996_));
 sky130_fd_sc_hd__clkbuf_1 _2174_ (.A(_0996_),
    .X(_0057_));
 sky130_fd_sc_hd__buf_4 _2175_ (.A(_0887_),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_1 _2176_ (.A0(_0997_),
    .A1(\RAM[14][2] ),
    .S(_0993_),
    .X(_0998_));
 sky130_fd_sc_hd__clkbuf_1 _2177_ (.A(_0998_),
    .X(_0058_));
 sky130_fd_sc_hd__clkbuf_4 _2178_ (.A(_0890_),
    .X(_0999_));
 sky130_fd_sc_hd__mux2_1 _2179_ (.A0(_0999_),
    .A1(\RAM[14][3] ),
    .S(_0993_),
    .X(_1000_));
 sky130_fd_sc_hd__clkbuf_1 _2180_ (.A(_1000_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _2181_ (.A(_0939_),
    .B(_0984_),
    .X(_1001_));
 sky130_fd_sc_hd__mux2_1 _2182_ (.A0(\RAM[15][0] ),
    .A1(_0876_),
    .S(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__clkbuf_1 _2183_ (.A(_1002_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _2184_ (.A0(\RAM[15][1] ),
    .A1(_0885_),
    .S(_1001_),
    .X(_1003_));
 sky130_fd_sc_hd__clkbuf_1 _2185_ (.A(_1003_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2186_ (.A0(\RAM[15][2] ),
    .A1(_0888_),
    .S(_1001_),
    .X(_1004_));
 sky130_fd_sc_hd__clkbuf_1 _2187_ (.A(_1004_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2188_ (.A0(\RAM[15][3] ),
    .A1(_0891_),
    .S(_1001_),
    .X(_1005_));
 sky130_fd_sc_hd__clkbuf_1 _2189_ (.A(_1005_),
    .X(_0063_));
 sky130_fd_sc_hd__or3_1 _2190_ (.A(_0539_),
    .B(_0558_),
    .C(_0556_),
    .X(_1006_));
 sky130_fd_sc_hd__buf_6 _2191_ (.A(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__nor2_2 _2192_ (.A(_0932_),
    .B(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__mux2_1 _2193_ (.A0(\RAM[16][0] ),
    .A1(_0876_),
    .S(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__clkbuf_1 _2194_ (.A(_1009_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _2195_ (.A0(\RAM[16][1] ),
    .A1(_0885_),
    .S(_1008_),
    .X(_1010_));
 sky130_fd_sc_hd__clkbuf_1 _2196_ (.A(_1010_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _2197_ (.A0(\RAM[16][2] ),
    .A1(_0888_),
    .S(_1008_),
    .X(_1011_));
 sky130_fd_sc_hd__clkbuf_1 _2198_ (.A(_1011_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _2199_ (.A0(\RAM[16][3] ),
    .A1(_0891_),
    .S(_1008_),
    .X(_1012_));
 sky130_fd_sc_hd__clkbuf_1 _2200_ (.A(_1012_),
    .X(_0067_));
 sky130_fd_sc_hd__nor2_2 _2201_ (.A(_0916_),
    .B(_0932_),
    .Y(_1013_));
 sky130_fd_sc_hd__mux2_1 _2202_ (.A0(\RAM[17][0] ),
    .A1(_0876_),
    .S(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__clkbuf_1 _2203_ (.A(_1014_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2204_ (.A0(\RAM[17][1] ),
    .A1(_0885_),
    .S(_1013_),
    .X(_1015_));
 sky130_fd_sc_hd__clkbuf_1 _2205_ (.A(_1015_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _2206_ (.A0(\RAM[17][2] ),
    .A1(_0888_),
    .S(_1013_),
    .X(_1016_));
 sky130_fd_sc_hd__clkbuf_1 _2207_ (.A(_1016_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _2208_ (.A0(\RAM[17][3] ),
    .A1(_0891_),
    .S(_1013_),
    .X(_1017_));
 sky130_fd_sc_hd__clkbuf_1 _2209_ (.A(_1017_),
    .X(_0071_));
 sky130_fd_sc_hd__clkbuf_4 _2210_ (.A(net8),
    .X(_1018_));
 sky130_fd_sc_hd__clkbuf_4 _2211_ (.A(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__or3_1 _2212_ (.A(_0539_),
    .B(_0524_),
    .C(_0556_),
    .X(_1020_));
 sky130_fd_sc_hd__buf_6 _2213_ (.A(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__nor2_2 _2214_ (.A(_0932_),
    .B(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__mux2_1 _2215_ (.A0(\RAM[18][0] ),
    .A1(_1019_),
    .S(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__clkbuf_1 _2216_ (.A(_1023_),
    .X(_0072_));
 sky130_fd_sc_hd__clkbuf_4 _2217_ (.A(net9),
    .X(_1024_));
 sky130_fd_sc_hd__buf_2 _2218_ (.A(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__mux2_1 _2219_ (.A0(\RAM[18][1] ),
    .A1(_1025_),
    .S(_1022_),
    .X(_1026_));
 sky130_fd_sc_hd__clkbuf_1 _2220_ (.A(_1026_),
    .X(_0073_));
 sky130_fd_sc_hd__clkbuf_4 _2221_ (.A(net10),
    .X(_1027_));
 sky130_fd_sc_hd__buf_2 _2222_ (.A(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__mux2_1 _2223_ (.A0(\RAM[18][2] ),
    .A1(_1028_),
    .S(_1022_),
    .X(_1029_));
 sky130_fd_sc_hd__clkbuf_1 _2224_ (.A(_1029_),
    .X(_0074_));
 sky130_fd_sc_hd__clkbuf_4 _2225_ (.A(net11),
    .X(_1030_));
 sky130_fd_sc_hd__buf_2 _2226_ (.A(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__mux2_1 _2227_ (.A0(\RAM[18][3] ),
    .A1(_1031_),
    .S(_1022_),
    .X(_1032_));
 sky130_fd_sc_hd__clkbuf_1 _2228_ (.A(_1032_),
    .X(_0075_));
 sky130_fd_sc_hd__nor2_2 _2229_ (.A(_0916_),
    .B(_0978_),
    .Y(_1033_));
 sky130_fd_sc_hd__mux2_1 _2230_ (.A0(\RAM[1][0] ),
    .A1(_1019_),
    .S(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__clkbuf_1 _2231_ (.A(_1034_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2232_ (.A0(\RAM[1][1] ),
    .A1(_1025_),
    .S(_1033_),
    .X(_1035_));
 sky130_fd_sc_hd__clkbuf_1 _2233_ (.A(_1035_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2234_ (.A0(\RAM[1][2] ),
    .A1(_1028_),
    .S(_1033_),
    .X(_1036_));
 sky130_fd_sc_hd__clkbuf_1 _2235_ (.A(_1036_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _2236_ (.A0(\RAM[1][3] ),
    .A1(_1031_),
    .S(_1033_),
    .X(_1037_));
 sky130_fd_sc_hd__clkbuf_1 _2237_ (.A(_1037_),
    .X(_0079_));
 sky130_fd_sc_hd__or3_1 _2238_ (.A(_0539_),
    .B(_0558_),
    .C(_0569_),
    .X(_1038_));
 sky130_fd_sc_hd__buf_6 _2239_ (.A(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__nor2_2 _2240_ (.A(_0932_),
    .B(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__mux2_1 _2241_ (.A0(\RAM[20][0] ),
    .A1(_1019_),
    .S(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__clkbuf_1 _2242_ (.A(_1041_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2243_ (.A0(\RAM[20][1] ),
    .A1(_1025_),
    .S(_1040_),
    .X(_1042_));
 sky130_fd_sc_hd__clkbuf_1 _2244_ (.A(_1042_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2245_ (.A0(\RAM[20][2] ),
    .A1(_1028_),
    .S(_1040_),
    .X(_1043_));
 sky130_fd_sc_hd__clkbuf_1 _2246_ (.A(_1043_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2247_ (.A0(\RAM[20][3] ),
    .A1(_1031_),
    .S(_1040_),
    .X(_1044_));
 sky130_fd_sc_hd__clkbuf_1 _2248_ (.A(_1044_),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_2 _2249_ (.A(_0878_),
    .B(_0932_),
    .Y(_1045_));
 sky130_fd_sc_hd__mux2_1 _2250_ (.A0(\RAM[21][0] ),
    .A1(_1019_),
    .S(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__clkbuf_1 _2251_ (.A(_1046_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2252_ (.A0(\RAM[21][1] ),
    .A1(_1025_),
    .S(_1045_),
    .X(_1047_));
 sky130_fd_sc_hd__clkbuf_1 _2253_ (.A(_1047_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2254_ (.A0(\RAM[21][2] ),
    .A1(_1028_),
    .S(_1045_),
    .X(_1048_));
 sky130_fd_sc_hd__clkbuf_1 _2255_ (.A(_1048_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2256_ (.A0(\RAM[21][3] ),
    .A1(_1031_),
    .S(_1045_),
    .X(_1049_));
 sky130_fd_sc_hd__clkbuf_1 _2257_ (.A(_1049_),
    .X(_0087_));
 sky130_fd_sc_hd__or3_1 _2258_ (.A(_0611_),
    .B(_0524_),
    .C(_0569_),
    .X(_1050_));
 sky130_fd_sc_hd__buf_4 _2259_ (.A(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__nor2_2 _2260_ (.A(_0932_),
    .B(_1051_),
    .Y(_1052_));
 sky130_fd_sc_hd__mux2_1 _2261_ (.A0(\RAM[22][0] ),
    .A1(_1019_),
    .S(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__clkbuf_1 _2262_ (.A(_1053_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2263_ (.A0(\RAM[22][1] ),
    .A1(_1025_),
    .S(_1052_),
    .X(_1054_));
 sky130_fd_sc_hd__clkbuf_1 _2264_ (.A(_1054_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2265_ (.A0(\RAM[22][2] ),
    .A1(_1028_),
    .S(_1052_),
    .X(_1055_));
 sky130_fd_sc_hd__clkbuf_1 _2266_ (.A(_1055_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _2267_ (.A0(\RAM[22][3] ),
    .A1(_1031_),
    .S(_1052_),
    .X(_1056_));
 sky130_fd_sc_hd__clkbuf_1 _2268_ (.A(_1056_),
    .X(_0091_));
 sky130_fd_sc_hd__nand2_2 _2269_ (.A(_0922_),
    .B(_0945_),
    .Y(_1057_));
 sky130_fd_sc_hd__mux2_1 _2270_ (.A0(_0990_),
    .A1(\RAM[23][0] ),
    .S(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__clkbuf_1 _2271_ (.A(_1058_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2272_ (.A0(_0995_),
    .A1(\RAM[23][1] ),
    .S(_1057_),
    .X(_1059_));
 sky130_fd_sc_hd__clkbuf_1 _2273_ (.A(_1059_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2274_ (.A0(_0997_),
    .A1(\RAM[23][2] ),
    .S(_1057_),
    .X(_1060_));
 sky130_fd_sc_hd__clkbuf_1 _2275_ (.A(_1060_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _2276_ (.A0(_0999_),
    .A1(\RAM[23][3] ),
    .S(_1057_),
    .X(_1061_));
 sky130_fd_sc_hd__clkbuf_1 _2277_ (.A(_1061_),
    .X(_0095_));
 sky130_fd_sc_hd__or3_1 _2278_ (.A(_0539_),
    .B(_0558_),
    .C(_0560_),
    .X(_1062_));
 sky130_fd_sc_hd__buf_8 _2279_ (.A(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__nor2_2 _2280_ (.A(_0932_),
    .B(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__mux2_1 _2281_ (.A0(\RAM[24][0] ),
    .A1(_1019_),
    .S(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__clkbuf_1 _2282_ (.A(_1065_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _2283_ (.A0(\RAM[24][1] ),
    .A1(_1025_),
    .S(_1064_),
    .X(_1066_));
 sky130_fd_sc_hd__clkbuf_1 _2284_ (.A(_1066_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _2285_ (.A0(\RAM[24][2] ),
    .A1(_1028_),
    .S(_1064_),
    .X(_1067_));
 sky130_fd_sc_hd__clkbuf_1 _2286_ (.A(_1067_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _2287_ (.A0(\RAM[24][3] ),
    .A1(_1031_),
    .S(_1064_),
    .X(_1068_));
 sky130_fd_sc_hd__clkbuf_1 _2288_ (.A(_1068_),
    .X(_0099_));
 sky130_fd_sc_hd__or2_4 _2289_ (.A(_0877_),
    .B(_0561_),
    .X(_1069_));
 sky130_fd_sc_hd__nor2_2 _2290_ (.A(_1069_),
    .B(_0932_),
    .Y(_1070_));
 sky130_fd_sc_hd__mux2_1 _2291_ (.A0(\RAM[25][0] ),
    .A1(_1019_),
    .S(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__clkbuf_1 _2292_ (.A(_1071_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2293_ (.A0(\RAM[25][1] ),
    .A1(_1025_),
    .S(_1070_),
    .X(_1072_));
 sky130_fd_sc_hd__clkbuf_1 _2294_ (.A(_1072_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2295_ (.A0(\RAM[25][2] ),
    .A1(_1028_),
    .S(_1070_),
    .X(_1073_));
 sky130_fd_sc_hd__clkbuf_1 _2296_ (.A(_1073_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _2297_ (.A0(\RAM[25][3] ),
    .A1(_1031_),
    .S(_1070_),
    .X(_1074_));
 sky130_fd_sc_hd__clkbuf_1 _2298_ (.A(_1074_),
    .X(_0103_));
 sky130_fd_sc_hd__or3_1 _2299_ (.A(_0611_),
    .B(_0524_),
    .C(_0560_),
    .X(_1075_));
 sky130_fd_sc_hd__buf_6 _2300_ (.A(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__nor2_2 _2301_ (.A(_0932_),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__mux2_1 _2302_ (.A0(\RAM[26][0] ),
    .A1(_1019_),
    .S(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__clkbuf_1 _2303_ (.A(_1078_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _2304_ (.A0(\RAM[26][1] ),
    .A1(_1025_),
    .S(_1077_),
    .X(_1079_));
 sky130_fd_sc_hd__clkbuf_1 _2305_ (.A(_1079_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2306_ (.A0(\RAM[26][2] ),
    .A1(_1028_),
    .S(_1077_),
    .X(_1080_));
 sky130_fd_sc_hd__clkbuf_1 _2307_ (.A(_1080_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _2308_ (.A0(\RAM[26][3] ),
    .A1(_1031_),
    .S(_1077_),
    .X(_1081_));
 sky130_fd_sc_hd__clkbuf_1 _2309_ (.A(_1081_),
    .X(_0107_));
 sky130_fd_sc_hd__nand2_2 _2310_ (.A(_0905_),
    .B(_0945_),
    .Y(_1082_));
 sky130_fd_sc_hd__mux2_1 _2311_ (.A0(_0990_),
    .A1(\RAM[27][0] ),
    .S(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__clkbuf_1 _2312_ (.A(_1083_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _2313_ (.A0(_0995_),
    .A1(\RAM[27][1] ),
    .S(_1082_),
    .X(_1084_));
 sky130_fd_sc_hd__clkbuf_1 _2314_ (.A(_1084_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _2315_ (.A0(_0997_),
    .A1(\RAM[27][2] ),
    .S(_1082_),
    .X(_1085_));
 sky130_fd_sc_hd__clkbuf_1 _2316_ (.A(_1085_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _2317_ (.A0(_0999_),
    .A1(\RAM[27][3] ),
    .S(_1082_),
    .X(_1086_));
 sky130_fd_sc_hd__clkbuf_1 _2318_ (.A(_1086_),
    .X(_0111_));
 sky130_fd_sc_hd__nor2_2 _2319_ (.A(_0931_),
    .B(_0976_),
    .Y(_1087_));
 sky130_fd_sc_hd__mux2_1 _2320_ (.A0(\RAM[28][0] ),
    .A1(_1019_),
    .S(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__clkbuf_1 _2321_ (.A(_1088_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _2322_ (.A0(\RAM[28][1] ),
    .A1(_1025_),
    .S(_1087_),
    .X(_1089_));
 sky130_fd_sc_hd__clkbuf_1 _2323_ (.A(_1089_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _2324_ (.A0(\RAM[28][2] ),
    .A1(_1028_),
    .S(_1087_),
    .X(_1090_));
 sky130_fd_sc_hd__clkbuf_1 _2325_ (.A(_1090_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _2326_ (.A0(\RAM[28][3] ),
    .A1(_1031_),
    .S(_1087_),
    .X(_1091_));
 sky130_fd_sc_hd__clkbuf_1 _2327_ (.A(_1091_),
    .X(_0115_));
 sky130_fd_sc_hd__nor2_2 _2328_ (.A(_0978_),
    .B(_1021_),
    .Y(_1092_));
 sky130_fd_sc_hd__mux2_1 _2329_ (.A0(\RAM[2][0] ),
    .A1(_1019_),
    .S(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__clkbuf_1 _2330_ (.A(_1093_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _2331_ (.A0(\RAM[2][1] ),
    .A1(_1025_),
    .S(_1092_),
    .X(_1094_));
 sky130_fd_sc_hd__clkbuf_1 _2332_ (.A(_1094_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _2333_ (.A0(\RAM[2][2] ),
    .A1(_1028_),
    .S(_1092_),
    .X(_1095_));
 sky130_fd_sc_hd__clkbuf_1 _2334_ (.A(_1095_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _2335_ (.A0(\RAM[2][3] ),
    .A1(_1031_),
    .S(_1092_),
    .X(_1096_));
 sky130_fd_sc_hd__clkbuf_1 _2336_ (.A(_1096_),
    .X(_0119_));
 sky130_fd_sc_hd__nand2_2 _2337_ (.A(_0945_),
    .B(_0992_),
    .Y(_1097_));
 sky130_fd_sc_hd__mux2_1 _2338_ (.A0(_0990_),
    .A1(\RAM[30][0] ),
    .S(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__clkbuf_1 _2339_ (.A(_1098_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _2340_ (.A0(_0995_),
    .A1(\RAM[30][1] ),
    .S(_1097_),
    .X(_1099_));
 sky130_fd_sc_hd__clkbuf_1 _2341_ (.A(_1099_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2342_ (.A0(_0997_),
    .A1(\RAM[30][2] ),
    .S(_1097_),
    .X(_1100_));
 sky130_fd_sc_hd__clkbuf_1 _2343_ (.A(_1100_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _2344_ (.A0(_0999_),
    .A1(\RAM[30][3] ),
    .S(_1097_),
    .X(_1101_));
 sky130_fd_sc_hd__clkbuf_1 _2345_ (.A(_1101_),
    .X(_0123_));
 sky130_fd_sc_hd__nand2_2 _2346_ (.A(_0945_),
    .B(_0939_),
    .Y(_1102_));
 sky130_fd_sc_hd__mux2_1 _2347_ (.A0(_0990_),
    .A1(\RAM[31][0] ),
    .S(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__clkbuf_1 _2348_ (.A(_1103_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _2349_ (.A0(_0995_),
    .A1(\RAM[31][1] ),
    .S(_1102_),
    .X(_1104_));
 sky130_fd_sc_hd__clkbuf_1 _2350_ (.A(_1104_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2351_ (.A0(_0997_),
    .A1(\RAM[31][2] ),
    .S(_1102_),
    .X(_1105_));
 sky130_fd_sc_hd__clkbuf_1 _2352_ (.A(_1105_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _2353_ (.A0(_0999_),
    .A1(\RAM[31][3] ),
    .S(_1102_),
    .X(_1106_));
 sky130_fd_sc_hd__clkbuf_1 _2354_ (.A(_1106_),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_4 _2355_ (.A(_1018_),
    .X(_1107_));
 sky130_fd_sc_hd__or2_1 _2356_ (.A(_0923_),
    .B(_0906_),
    .X(_1108_));
 sky130_fd_sc_hd__buf_4 _2357_ (.A(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__nor2_2 _2358_ (.A(_1109_),
    .B(_1007_),
    .Y(_1110_));
 sky130_fd_sc_hd__mux2_1 _2359_ (.A0(\RAM[32][0] ),
    .A1(_1107_),
    .S(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__clkbuf_1 _2360_ (.A(_1111_),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_4 _2361_ (.A(_1024_),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_1 _2362_ (.A0(\RAM[32][1] ),
    .A1(_1112_),
    .S(_1110_),
    .X(_1113_));
 sky130_fd_sc_hd__clkbuf_1 _2363_ (.A(_1113_),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_4 _2364_ (.A(_1027_),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_1 _2365_ (.A0(\RAM[32][2] ),
    .A1(_1114_),
    .S(_1110_),
    .X(_1115_));
 sky130_fd_sc_hd__clkbuf_1 _2366_ (.A(_1115_),
    .X(_0130_));
 sky130_fd_sc_hd__buf_2 _2367_ (.A(_1030_),
    .X(_1116_));
 sky130_fd_sc_hd__mux2_1 _2368_ (.A0(\RAM[32][3] ),
    .A1(_1116_),
    .S(_1110_),
    .X(_1117_));
 sky130_fd_sc_hd__clkbuf_1 _2369_ (.A(_1117_),
    .X(_0131_));
 sky130_fd_sc_hd__nor2_2 _2370_ (.A(_0916_),
    .B(_1109_),
    .Y(_1118_));
 sky130_fd_sc_hd__mux2_1 _2371_ (.A0(\RAM[33][0] ),
    .A1(_1107_),
    .S(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__clkbuf_1 _2372_ (.A(_1119_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2373_ (.A0(\RAM[33][1] ),
    .A1(_1112_),
    .S(_1118_),
    .X(_1120_));
 sky130_fd_sc_hd__clkbuf_1 _2374_ (.A(_1120_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _2375_ (.A0(\RAM[33][2] ),
    .A1(_1114_),
    .S(_1118_),
    .X(_1121_));
 sky130_fd_sc_hd__clkbuf_1 _2376_ (.A(_1121_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _2377_ (.A0(\RAM[33][3] ),
    .A1(_1116_),
    .S(_1118_),
    .X(_1122_));
 sky130_fd_sc_hd__clkbuf_1 _2378_ (.A(_1122_),
    .X(_0135_));
 sky130_fd_sc_hd__nor2_2 _2379_ (.A(_1109_),
    .B(_1021_),
    .Y(_1123_));
 sky130_fd_sc_hd__mux2_1 _2380_ (.A0(\RAM[34][0] ),
    .A1(_1107_),
    .S(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__clkbuf_1 _2381_ (.A(_1124_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _2382_ (.A0(\RAM[34][1] ),
    .A1(_1112_),
    .S(_1123_),
    .X(_1125_));
 sky130_fd_sc_hd__clkbuf_1 _2383_ (.A(_1125_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _2384_ (.A0(\RAM[34][2] ),
    .A1(_1114_),
    .S(_1123_),
    .X(_1126_));
 sky130_fd_sc_hd__clkbuf_1 _2385_ (.A(_1126_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _2386_ (.A0(\RAM[34][3] ),
    .A1(_1116_),
    .S(_1123_),
    .X(_1127_));
 sky130_fd_sc_hd__clkbuf_1 _2387_ (.A(_1127_),
    .X(_0139_));
 sky130_fd_sc_hd__nor2_2 _2388_ (.A(_1109_),
    .B(_0930_),
    .Y(_1128_));
 sky130_fd_sc_hd__mux2_1 _2389_ (.A0(\RAM[35][0] ),
    .A1(_1107_),
    .S(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__clkbuf_1 _2390_ (.A(_1129_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _2391_ (.A0(\RAM[35][1] ),
    .A1(_1112_),
    .S(_1128_),
    .X(_1130_));
 sky130_fd_sc_hd__clkbuf_1 _2392_ (.A(_1130_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2393_ (.A0(\RAM[35][2] ),
    .A1(_1114_),
    .S(_1128_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_1 _2394_ (.A(_1131_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _2395_ (.A0(\RAM[35][3] ),
    .A1(_1116_),
    .S(_1128_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _2396_ (.A(_1132_),
    .X(_0143_));
 sky130_fd_sc_hd__nor2_2 _2397_ (.A(_1109_),
    .B(_1039_),
    .Y(_1133_));
 sky130_fd_sc_hd__mux2_1 _2398_ (.A0(\RAM[36][0] ),
    .A1(_1107_),
    .S(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _2399_ (.A(_1134_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2400_ (.A0(\RAM[36][1] ),
    .A1(_1112_),
    .S(_1133_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_1 _2401_ (.A(_1135_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2402_ (.A0(\RAM[36][2] ),
    .A1(_1114_),
    .S(_1133_),
    .X(_1136_));
 sky130_fd_sc_hd__clkbuf_1 _2403_ (.A(_1136_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2404_ (.A0(\RAM[36][3] ),
    .A1(_1116_),
    .S(_1133_),
    .X(_1137_));
 sky130_fd_sc_hd__clkbuf_1 _2405_ (.A(_1137_),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_2 _2406_ (.A(_0878_),
    .B(_1109_),
    .Y(_1138_));
 sky130_fd_sc_hd__mux2_1 _2407_ (.A0(\RAM[37][0] ),
    .A1(_1107_),
    .S(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__clkbuf_1 _2408_ (.A(_1139_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2409_ (.A0(\RAM[37][1] ),
    .A1(_1112_),
    .S(_1138_),
    .X(_1140_));
 sky130_fd_sc_hd__clkbuf_1 _2410_ (.A(_1140_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(\RAM[37][2] ),
    .A1(_1114_),
    .S(_1138_),
    .X(_1141_));
 sky130_fd_sc_hd__clkbuf_1 _2412_ (.A(_1141_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2413_ (.A0(\RAM[37][3] ),
    .A1(_1116_),
    .S(_1138_),
    .X(_1142_));
 sky130_fd_sc_hd__clkbuf_1 _2414_ (.A(_1142_),
    .X(_0151_));
 sky130_fd_sc_hd__nor2_2 _2415_ (.A(_1109_),
    .B(_1051_),
    .Y(_1143_));
 sky130_fd_sc_hd__mux2_1 _2416_ (.A0(\RAM[38][0] ),
    .A1(_1107_),
    .S(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__clkbuf_1 _2417_ (.A(_1144_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2418_ (.A0(\RAM[38][1] ),
    .A1(_1112_),
    .S(_1143_),
    .X(_1145_));
 sky130_fd_sc_hd__clkbuf_1 _2419_ (.A(_1145_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2420_ (.A0(\RAM[38][2] ),
    .A1(_1114_),
    .S(_1143_),
    .X(_1146_));
 sky130_fd_sc_hd__clkbuf_1 _2421_ (.A(_1146_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2422_ (.A0(\RAM[38][3] ),
    .A1(_1116_),
    .S(_1143_),
    .X(_1147_));
 sky130_fd_sc_hd__clkbuf_1 _2423_ (.A(_1147_),
    .X(_0155_));
 sky130_fd_sc_hd__nor2_2 _2424_ (.A(_0930_),
    .B(_0978_),
    .Y(_1148_));
 sky130_fd_sc_hd__mux2_1 _2425_ (.A0(\RAM[3][0] ),
    .A1(_1107_),
    .S(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__clkbuf_1 _2426_ (.A(_1149_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2427_ (.A0(\RAM[3][1] ),
    .A1(_1112_),
    .S(_1148_),
    .X(_1150_));
 sky130_fd_sc_hd__clkbuf_1 _2428_ (.A(_1150_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2429_ (.A0(\RAM[3][2] ),
    .A1(_1114_),
    .S(_1148_),
    .X(_1151_));
 sky130_fd_sc_hd__clkbuf_1 _2430_ (.A(_1151_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2431_ (.A0(\RAM[3][3] ),
    .A1(_1116_),
    .S(_1148_),
    .X(_1152_));
 sky130_fd_sc_hd__clkbuf_1 _2432_ (.A(_1152_),
    .X(_0159_));
 sky130_fd_sc_hd__nor2_2 _2433_ (.A(_1109_),
    .B(_1063_),
    .Y(_1153_));
 sky130_fd_sc_hd__mux2_1 _2434_ (.A0(\RAM[40][0] ),
    .A1(_1107_),
    .S(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__clkbuf_1 _2435_ (.A(_1154_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2436_ (.A0(\RAM[40][1] ),
    .A1(_1112_),
    .S(_1153_),
    .X(_1155_));
 sky130_fd_sc_hd__clkbuf_1 _2437_ (.A(_1155_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(\RAM[40][2] ),
    .A1(_1114_),
    .S(_1153_),
    .X(_1156_));
 sky130_fd_sc_hd__clkbuf_1 _2439_ (.A(_1156_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2440_ (.A0(\RAM[40][3] ),
    .A1(_1116_),
    .S(_1153_),
    .X(_1157_));
 sky130_fd_sc_hd__clkbuf_1 _2441_ (.A(_1157_),
    .X(_0163_));
 sky130_fd_sc_hd__nor2_2 _2442_ (.A(_1069_),
    .B(_1109_),
    .Y(_1158_));
 sky130_fd_sc_hd__mux2_1 _2443_ (.A0(\RAM[41][0] ),
    .A1(_1107_),
    .S(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__clkbuf_1 _2444_ (.A(_1159_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2445_ (.A0(\RAM[41][1] ),
    .A1(_1112_),
    .S(_1158_),
    .X(_1160_));
 sky130_fd_sc_hd__clkbuf_1 _2446_ (.A(_1160_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _2447_ (.A0(\RAM[41][2] ),
    .A1(_1114_),
    .S(_1158_),
    .X(_1161_));
 sky130_fd_sc_hd__clkbuf_1 _2448_ (.A(_1161_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2449_ (.A0(\RAM[41][3] ),
    .A1(_1116_),
    .S(_1158_),
    .X(_1162_));
 sky130_fd_sc_hd__clkbuf_1 _2450_ (.A(_1162_),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_4 _2451_ (.A(_0875_),
    .X(_1163_));
 sky130_fd_sc_hd__nor2_2 _2452_ (.A(_1109_),
    .B(_1076_),
    .Y(_1164_));
 sky130_fd_sc_hd__mux2_1 _2453_ (.A0(\RAM[42][0] ),
    .A1(_1163_),
    .S(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__clkbuf_1 _2454_ (.A(_1165_),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_4 _2455_ (.A(_0884_),
    .X(_1166_));
 sky130_fd_sc_hd__mux2_1 _2456_ (.A0(\RAM[42][1] ),
    .A1(_1166_),
    .S(_1164_),
    .X(_1167_));
 sky130_fd_sc_hd__clkbuf_1 _2457_ (.A(_1167_),
    .X(_0169_));
 sky130_fd_sc_hd__clkbuf_4 _2458_ (.A(_0887_),
    .X(_1168_));
 sky130_fd_sc_hd__mux2_1 _2459_ (.A0(\RAM[42][2] ),
    .A1(_1168_),
    .S(_1164_),
    .X(_1169_));
 sky130_fd_sc_hd__clkbuf_1 _2460_ (.A(_1169_),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_4 _2461_ (.A(_0890_),
    .X(_1170_));
 sky130_fd_sc_hd__mux2_1 _2462_ (.A0(\RAM[42][3] ),
    .A1(_1170_),
    .S(_1164_),
    .X(_1171_));
 sky130_fd_sc_hd__clkbuf_1 _2463_ (.A(_1171_),
    .X(_0171_));
 sky130_fd_sc_hd__nand2_2 _2464_ (.A(_0905_),
    .B(_0924_),
    .Y(_1172_));
 sky130_fd_sc_hd__mux2_1 _2465_ (.A0(_0990_),
    .A1(\RAM[43][0] ),
    .S(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_1 _2466_ (.A(_1173_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2467_ (.A0(_0995_),
    .A1(\RAM[43][1] ),
    .S(_1172_),
    .X(_1174_));
 sky130_fd_sc_hd__clkbuf_1 _2468_ (.A(_1174_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2469_ (.A0(_0997_),
    .A1(\RAM[43][2] ),
    .S(_1172_),
    .X(_1175_));
 sky130_fd_sc_hd__clkbuf_1 _2470_ (.A(_1175_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _2471_ (.A0(_0999_),
    .A1(\RAM[43][3] ),
    .S(_1172_),
    .X(_1176_));
 sky130_fd_sc_hd__clkbuf_1 _2472_ (.A(_1176_),
    .X(_0175_));
 sky130_fd_sc_hd__nor2_2 _2473_ (.A(_1108_),
    .B(_0976_),
    .Y(_1177_));
 sky130_fd_sc_hd__mux2_1 _2474_ (.A0(\RAM[44][0] ),
    .A1(_1163_),
    .S(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__clkbuf_1 _2475_ (.A(_1178_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2476_ (.A0(\RAM[44][1] ),
    .A1(_1166_),
    .S(_1177_),
    .X(_1179_));
 sky130_fd_sc_hd__clkbuf_1 _2477_ (.A(_1179_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2478_ (.A0(\RAM[44][2] ),
    .A1(_1168_),
    .S(_1177_),
    .X(_1180_));
 sky130_fd_sc_hd__clkbuf_1 _2479_ (.A(_1180_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2480_ (.A0(\RAM[44][3] ),
    .A1(_1170_),
    .S(_1177_),
    .X(_1181_));
 sky130_fd_sc_hd__clkbuf_1 _2481_ (.A(_1181_),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_2 _2482_ (.A(_0924_),
    .B(_0946_),
    .Y(_1182_));
 sky130_fd_sc_hd__mux2_1 _2483_ (.A0(_0990_),
    .A1(\RAM[45][0] ),
    .S(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__clkbuf_1 _2484_ (.A(_1183_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2485_ (.A0(_0995_),
    .A1(\RAM[45][1] ),
    .S(_1182_),
    .X(_1184_));
 sky130_fd_sc_hd__clkbuf_1 _2486_ (.A(_1184_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _2487_ (.A0(_0997_),
    .A1(\RAM[45][2] ),
    .S(_1182_),
    .X(_1185_));
 sky130_fd_sc_hd__clkbuf_1 _2488_ (.A(_1185_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2489_ (.A0(_0999_),
    .A1(\RAM[45][3] ),
    .S(_1182_),
    .X(_1186_));
 sky130_fd_sc_hd__clkbuf_1 _2490_ (.A(_1186_),
    .X(_0183_));
 sky130_fd_sc_hd__nand2_2 _2491_ (.A(_0924_),
    .B(_0992_),
    .Y(_1187_));
 sky130_fd_sc_hd__mux2_1 _2492_ (.A0(_0990_),
    .A1(\RAM[46][0] ),
    .S(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__clkbuf_1 _2493_ (.A(_1188_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _2494_ (.A0(_0995_),
    .A1(\RAM[46][1] ),
    .S(_1187_),
    .X(_1189_));
 sky130_fd_sc_hd__clkbuf_1 _2495_ (.A(_1189_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _2496_ (.A0(_0997_),
    .A1(\RAM[46][2] ),
    .S(_1187_),
    .X(_1190_));
 sky130_fd_sc_hd__clkbuf_1 _2497_ (.A(_1190_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2498_ (.A0(_0999_),
    .A1(\RAM[46][3] ),
    .S(_1187_),
    .X(_1191_));
 sky130_fd_sc_hd__clkbuf_1 _2499_ (.A(_1191_),
    .X(_0187_));
 sky130_fd_sc_hd__nand2_2 _2500_ (.A(_0924_),
    .B(_0939_),
    .Y(_1192_));
 sky130_fd_sc_hd__mux2_1 _2501_ (.A0(_0990_),
    .A1(\RAM[47][0] ),
    .S(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__clkbuf_1 _2502_ (.A(_1193_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _2503_ (.A0(_0995_),
    .A1(\RAM[47][1] ),
    .S(_1192_),
    .X(_1194_));
 sky130_fd_sc_hd__clkbuf_1 _2504_ (.A(_1194_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _2505_ (.A0(_0997_),
    .A1(\RAM[47][2] ),
    .S(_1192_),
    .X(_1195_));
 sky130_fd_sc_hd__clkbuf_1 _2506_ (.A(_1195_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _2507_ (.A0(_0999_),
    .A1(\RAM[47][3] ),
    .S(_1192_),
    .X(_1196_));
 sky130_fd_sc_hd__clkbuf_1 _2508_ (.A(_1196_),
    .X(_0191_));
 sky130_fd_sc_hd__nor2_2 _2509_ (.A(_0914_),
    .B(_1007_),
    .Y(_1197_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(\RAM[48][0] ),
    .A1(_1163_),
    .S(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__clkbuf_1 _2511_ (.A(_1198_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(\RAM[48][1] ),
    .A1(_1166_),
    .S(_1197_),
    .X(_1199_));
 sky130_fd_sc_hd__clkbuf_1 _2513_ (.A(_1199_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _2514_ (.A0(\RAM[48][2] ),
    .A1(_1168_),
    .S(_1197_),
    .X(_1200_));
 sky130_fd_sc_hd__clkbuf_1 _2515_ (.A(_1200_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _2516_ (.A0(\RAM[48][3] ),
    .A1(_1170_),
    .S(_1197_),
    .X(_1201_));
 sky130_fd_sc_hd__clkbuf_1 _2517_ (.A(_1201_),
    .X(_0195_));
 sky130_fd_sc_hd__nor2_2 _2518_ (.A(_0978_),
    .B(_1039_),
    .Y(_1202_));
 sky130_fd_sc_hd__mux2_1 _2519_ (.A0(\RAM[4][0] ),
    .A1(_1163_),
    .S(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__clkbuf_1 _2520_ (.A(_1203_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _2521_ (.A0(\RAM[4][1] ),
    .A1(_1166_),
    .S(_1202_),
    .X(_1204_));
 sky130_fd_sc_hd__clkbuf_1 _2522_ (.A(_1204_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(\RAM[4][2] ),
    .A1(_1168_),
    .S(_1202_),
    .X(_1205_));
 sky130_fd_sc_hd__clkbuf_1 _2524_ (.A(_1205_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(\RAM[4][3] ),
    .A1(_1170_),
    .S(_1202_),
    .X(_1206_));
 sky130_fd_sc_hd__clkbuf_1 _2526_ (.A(_1206_),
    .X(_0199_));
 sky130_fd_sc_hd__nor2_2 _2527_ (.A(_0914_),
    .B(_1021_),
    .Y(_1207_));
 sky130_fd_sc_hd__mux2_1 _2528_ (.A0(\RAM[50][0] ),
    .A1(_1163_),
    .S(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__clkbuf_1 _2529_ (.A(_1208_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(\RAM[50][1] ),
    .A1(_1166_),
    .S(_1207_),
    .X(_1209_));
 sky130_fd_sc_hd__clkbuf_1 _2531_ (.A(_1209_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2532_ (.A0(\RAM[50][2] ),
    .A1(_1168_),
    .S(_1207_),
    .X(_1210_));
 sky130_fd_sc_hd__clkbuf_1 _2533_ (.A(_1210_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _2534_ (.A0(\RAM[50][3] ),
    .A1(_1170_),
    .S(_1207_),
    .X(_1211_));
 sky130_fd_sc_hd__clkbuf_1 _2535_ (.A(_1211_),
    .X(_0203_));
 sky130_fd_sc_hd__nand2_2 _2536_ (.A(_0907_),
    .B(_0952_),
    .Y(_1212_));
 sky130_fd_sc_hd__mux2_1 _2537_ (.A0(_0990_),
    .A1(\RAM[51][0] ),
    .S(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__clkbuf_1 _2538_ (.A(_1213_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _2539_ (.A0(_0995_),
    .A1(\RAM[51][1] ),
    .S(_1212_),
    .X(_1214_));
 sky130_fd_sc_hd__clkbuf_1 _2540_ (.A(_1214_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _2541_ (.A0(_0997_),
    .A1(\RAM[51][2] ),
    .S(_1212_),
    .X(_1215_));
 sky130_fd_sc_hd__clkbuf_1 _2542_ (.A(_1215_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _2543_ (.A0(_0999_),
    .A1(\RAM[51][3] ),
    .S(_1212_),
    .X(_1216_));
 sky130_fd_sc_hd__clkbuf_1 _2544_ (.A(_1216_),
    .X(_0207_));
 sky130_fd_sc_hd__nor2_2 _2545_ (.A(_0914_),
    .B(_1039_),
    .Y(_1217_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(\RAM[52][0] ),
    .A1(_1163_),
    .S(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__clkbuf_1 _2547_ (.A(_1218_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(\RAM[52][1] ),
    .A1(_1166_),
    .S(_1217_),
    .X(_1219_));
 sky130_fd_sc_hd__clkbuf_1 _2549_ (.A(_1219_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(\RAM[52][2] ),
    .A1(_1168_),
    .S(_1217_),
    .X(_1220_));
 sky130_fd_sc_hd__clkbuf_1 _2551_ (.A(_1220_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _2552_ (.A0(\RAM[52][3] ),
    .A1(_1170_),
    .S(_1217_),
    .X(_1221_));
 sky130_fd_sc_hd__clkbuf_1 _2553_ (.A(_1221_),
    .X(_0211_));
 sky130_fd_sc_hd__buf_2 _2554_ (.A(_0875_),
    .X(_1222_));
 sky130_fd_sc_hd__nor2_4 _2555_ (.A(_0570_),
    .B(_0877_),
    .Y(_1223_));
 sky130_fd_sc_hd__nand2_2 _2556_ (.A(_1223_),
    .B(_0907_),
    .Y(_1224_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(_1222_),
    .A1(\RAM[53][0] ),
    .S(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__clkbuf_1 _2558_ (.A(_1225_),
    .X(_0212_));
 sky130_fd_sc_hd__buf_2 _2559_ (.A(_0884_),
    .X(_1226_));
 sky130_fd_sc_hd__mux2_1 _2560_ (.A0(_1226_),
    .A1(\RAM[53][1] ),
    .S(_1224_),
    .X(_1227_));
 sky130_fd_sc_hd__clkbuf_1 _2561_ (.A(_1227_),
    .X(_0213_));
 sky130_fd_sc_hd__buf_2 _2562_ (.A(_0887_),
    .X(_1228_));
 sky130_fd_sc_hd__mux2_1 _2563_ (.A0(_1228_),
    .A1(\RAM[53][2] ),
    .S(_1224_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _2564_ (.A(_1229_),
    .X(_0214_));
 sky130_fd_sc_hd__buf_2 _2565_ (.A(_0890_),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_1 _2566_ (.A0(_1230_),
    .A1(\RAM[53][3] ),
    .S(_1224_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _2567_ (.A(_1231_),
    .X(_0215_));
 sky130_fd_sc_hd__or2_2 _2568_ (.A(_0914_),
    .B(_1051_),
    .X(_1232_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(_1222_),
    .A1(\RAM[54][0] ),
    .S(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__clkbuf_1 _2570_ (.A(_1233_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _2571_ (.A0(_1226_),
    .A1(\RAM[54][1] ),
    .S(_1232_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _2572_ (.A(_1234_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(_1228_),
    .A1(\RAM[54][2] ),
    .S(_1232_),
    .X(_1235_));
 sky130_fd_sc_hd__clkbuf_1 _2574_ (.A(_1235_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _2575_ (.A0(_1230_),
    .A1(\RAM[54][3] ),
    .S(_1232_),
    .X(_1236_));
 sky130_fd_sc_hd__clkbuf_1 _2576_ (.A(_1236_),
    .X(_0219_));
 sky130_fd_sc_hd__nand2_2 _2577_ (.A(_0907_),
    .B(_0922_),
    .Y(_1237_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(_1222_),
    .A1(\RAM[55][0] ),
    .S(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__clkbuf_1 _2579_ (.A(_1238_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(_1226_),
    .A1(\RAM[55][1] ),
    .S(_1237_),
    .X(_1239_));
 sky130_fd_sc_hd__clkbuf_1 _2581_ (.A(_1239_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(_1228_),
    .A1(\RAM[55][2] ),
    .S(_1237_),
    .X(_1240_));
 sky130_fd_sc_hd__clkbuf_1 _2583_ (.A(_1240_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _2584_ (.A0(_1230_),
    .A1(\RAM[55][3] ),
    .S(_1237_),
    .X(_1241_));
 sky130_fd_sc_hd__clkbuf_1 _2585_ (.A(_1241_),
    .X(_0223_));
 sky130_fd_sc_hd__nor2_2 _2586_ (.A(_0914_),
    .B(_1063_),
    .Y(_1242_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(\RAM[56][0] ),
    .A1(_1163_),
    .S(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__clkbuf_1 _2588_ (.A(_1243_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _2589_ (.A0(\RAM[56][1] ),
    .A1(_1166_),
    .S(_1242_),
    .X(_1244_));
 sky130_fd_sc_hd__clkbuf_1 _2590_ (.A(_1244_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _2591_ (.A0(\RAM[56][2] ),
    .A1(_1168_),
    .S(_1242_),
    .X(_1245_));
 sky130_fd_sc_hd__clkbuf_1 _2592_ (.A(_1245_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _2593_ (.A0(\RAM[56][3] ),
    .A1(_1170_),
    .S(_1242_),
    .X(_1246_));
 sky130_fd_sc_hd__clkbuf_1 _2594_ (.A(_1246_),
    .X(_0227_));
 sky130_fd_sc_hd__nand2_2 _2595_ (.A(_0894_),
    .B(_0907_),
    .Y(_1247_));
 sky130_fd_sc_hd__mux2_1 _2596_ (.A0(_1222_),
    .A1(\RAM[57][0] ),
    .S(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__clkbuf_1 _2597_ (.A(_1248_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _2598_ (.A0(_1226_),
    .A1(\RAM[57][1] ),
    .S(_1247_),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_1 _2599_ (.A(_1249_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _2600_ (.A0(_1228_),
    .A1(\RAM[57][2] ),
    .S(_1247_),
    .X(_1250_));
 sky130_fd_sc_hd__clkbuf_1 _2601_ (.A(_1250_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _2602_ (.A0(_1230_),
    .A1(\RAM[57][3] ),
    .S(_1247_),
    .X(_1251_));
 sky130_fd_sc_hd__clkbuf_1 _2603_ (.A(_1251_),
    .X(_0231_));
 sky130_fd_sc_hd__or2_2 _2604_ (.A(_0914_),
    .B(_1076_),
    .X(_1252_));
 sky130_fd_sc_hd__mux2_1 _2605_ (.A0(_1222_),
    .A1(\RAM[58][0] ),
    .S(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__clkbuf_1 _2606_ (.A(_1253_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _2607_ (.A0(_1226_),
    .A1(\RAM[58][1] ),
    .S(_1252_),
    .X(_1254_));
 sky130_fd_sc_hd__clkbuf_1 _2608_ (.A(_1254_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(_1228_),
    .A1(\RAM[58][2] ),
    .S(_1252_),
    .X(_1255_));
 sky130_fd_sc_hd__clkbuf_1 _2610_ (.A(_1255_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(_1230_),
    .A1(\RAM[58][3] ),
    .S(_1252_),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_1 _2612_ (.A(_1256_),
    .X(_0235_));
 sky130_fd_sc_hd__nor2_2 _2613_ (.A(_0878_),
    .B(_0978_),
    .Y(_1257_));
 sky130_fd_sc_hd__mux2_1 _2614_ (.A0(\RAM[5][0] ),
    .A1(_1163_),
    .S(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__clkbuf_1 _2615_ (.A(_1258_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _2616_ (.A0(\RAM[5][1] ),
    .A1(_1166_),
    .S(_1257_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_1 _2617_ (.A(_1259_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _2618_ (.A0(\RAM[5][2] ),
    .A1(_1168_),
    .S(_1257_),
    .X(_1260_));
 sky130_fd_sc_hd__clkbuf_1 _2619_ (.A(_1260_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _2620_ (.A0(\RAM[5][3] ),
    .A1(_1170_),
    .S(_1257_),
    .X(_1261_));
 sky130_fd_sc_hd__clkbuf_1 _2621_ (.A(_1261_),
    .X(_0239_));
 sky130_fd_sc_hd__or2_2 _2622_ (.A(_0914_),
    .B(_0976_),
    .X(_1262_));
 sky130_fd_sc_hd__mux2_1 _2623_ (.A0(_1222_),
    .A1(\RAM[60][0] ),
    .S(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__clkbuf_1 _2624_ (.A(_1263_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2625_ (.A0(_1226_),
    .A1(\RAM[60][1] ),
    .S(_1262_),
    .X(_1264_));
 sky130_fd_sc_hd__clkbuf_1 _2626_ (.A(_1264_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _2627_ (.A0(_1228_),
    .A1(\RAM[60][2] ),
    .S(_1262_),
    .X(_1265_));
 sky130_fd_sc_hd__clkbuf_1 _2628_ (.A(_1265_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _2629_ (.A0(_1230_),
    .A1(\RAM[60][3] ),
    .S(_1262_),
    .X(_1266_));
 sky130_fd_sc_hd__clkbuf_1 _2630_ (.A(_1266_),
    .X(_0243_));
 sky130_fd_sc_hd__nand2_2 _2631_ (.A(_0907_),
    .B(_0946_),
    .Y(_1267_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(_1222_),
    .A1(\RAM[61][0] ),
    .S(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_1 _2633_ (.A(_1268_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(_1226_),
    .A1(\RAM[61][1] ),
    .S(_1267_),
    .X(_1269_));
 sky130_fd_sc_hd__clkbuf_1 _2635_ (.A(_1269_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(_1228_),
    .A1(\RAM[61][2] ),
    .S(_1267_),
    .X(_1270_));
 sky130_fd_sc_hd__clkbuf_1 _2637_ (.A(_1270_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _2638_ (.A0(_1230_),
    .A1(\RAM[61][3] ),
    .S(_1267_),
    .X(_1271_));
 sky130_fd_sc_hd__clkbuf_1 _2639_ (.A(_1271_),
    .X(_0247_));
 sky130_fd_sc_hd__nand2_2 _2640_ (.A(_0907_),
    .B(_0992_),
    .Y(_1272_));
 sky130_fd_sc_hd__mux2_1 _2641_ (.A0(_1222_),
    .A1(\RAM[62][0] ),
    .S(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__clkbuf_1 _2642_ (.A(_1273_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _2643_ (.A0(_1226_),
    .A1(\RAM[62][1] ),
    .S(_1272_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _2644_ (.A(_1274_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(_1228_),
    .A1(\RAM[62][2] ),
    .S(_1272_),
    .X(_1275_));
 sky130_fd_sc_hd__clkbuf_1 _2646_ (.A(_1275_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _2647_ (.A0(_1230_),
    .A1(\RAM[62][3] ),
    .S(_1272_),
    .X(_1276_));
 sky130_fd_sc_hd__clkbuf_1 _2648_ (.A(_1276_),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_2 _2649_ (.A(_0907_),
    .B(_0939_),
    .Y(_1277_));
 sky130_fd_sc_hd__mux2_1 _2650_ (.A0(_1222_),
    .A1(\RAM[63][0] ),
    .S(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__clkbuf_1 _2651_ (.A(_1278_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _2652_ (.A0(_1226_),
    .A1(\RAM[63][1] ),
    .S(_1277_),
    .X(_1279_));
 sky130_fd_sc_hd__clkbuf_1 _2653_ (.A(_1279_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _2654_ (.A0(_1228_),
    .A1(\RAM[63][2] ),
    .S(_1277_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _2655_ (.A(_1280_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _2656_ (.A0(_1230_),
    .A1(\RAM[63][3] ),
    .S(_1277_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_1 _2657_ (.A(_1281_),
    .X(_0255_));
 sky130_fd_sc_hd__nor2_2 _2658_ (.A(_0881_),
    .B(_1007_),
    .Y(_1282_));
 sky130_fd_sc_hd__mux2_1 _2659_ (.A0(\RAM[64][0] ),
    .A1(_1163_),
    .S(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__clkbuf_1 _2660_ (.A(_1283_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _2661_ (.A0(\RAM[64][1] ),
    .A1(_1166_),
    .S(_1282_),
    .X(_1284_));
 sky130_fd_sc_hd__clkbuf_1 _2662_ (.A(_1284_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _2663_ (.A0(\RAM[64][2] ),
    .A1(_1168_),
    .S(_1282_),
    .X(_1285_));
 sky130_fd_sc_hd__clkbuf_1 _2664_ (.A(_1285_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _2665_ (.A0(\RAM[64][3] ),
    .A1(_1170_),
    .S(_1282_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_1 _2666_ (.A(_1286_),
    .X(_0259_));
 sky130_fd_sc_hd__nor2_2 _2667_ (.A(_0881_),
    .B(_0916_),
    .Y(_1287_));
 sky130_fd_sc_hd__mux2_1 _2668_ (.A0(\RAM[65][0] ),
    .A1(_1163_),
    .S(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_1 _2669_ (.A(_1288_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _2670_ (.A0(\RAM[65][1] ),
    .A1(_1166_),
    .S(_1287_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _2671_ (.A(_1289_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _2672_ (.A0(\RAM[65][2] ),
    .A1(_1168_),
    .S(_1287_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _2673_ (.A(_1290_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _2674_ (.A0(\RAM[65][3] ),
    .A1(_1170_),
    .S(_1287_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _2675_ (.A(_1291_),
    .X(_0263_));
 sky130_fd_sc_hd__clkbuf_4 _2676_ (.A(_0875_),
    .X(_1292_));
 sky130_fd_sc_hd__nor2_2 _2677_ (.A(_0881_),
    .B(_1021_),
    .Y(_1293_));
 sky130_fd_sc_hd__mux2_1 _2678_ (.A0(\RAM[66][0] ),
    .A1(_1292_),
    .S(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _2679_ (.A(_1294_),
    .X(_0264_));
 sky130_fd_sc_hd__clkbuf_4 _2680_ (.A(_0884_),
    .X(_1295_));
 sky130_fd_sc_hd__mux2_1 _2681_ (.A0(\RAM[66][1] ),
    .A1(_1295_),
    .S(_1293_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _2682_ (.A(_1296_),
    .X(_0265_));
 sky130_fd_sc_hd__clkbuf_4 _2683_ (.A(_0887_),
    .X(_1297_));
 sky130_fd_sc_hd__mux2_1 _2684_ (.A0(\RAM[66][2] ),
    .A1(_1297_),
    .S(_1293_),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_1 _2685_ (.A(_1298_),
    .X(_0266_));
 sky130_fd_sc_hd__clkbuf_4 _2686_ (.A(_0890_),
    .X(_1299_));
 sky130_fd_sc_hd__mux2_1 _2687_ (.A0(\RAM[66][3] ),
    .A1(_1299_),
    .S(_1293_),
    .X(_1300_));
 sky130_fd_sc_hd__clkbuf_1 _2688_ (.A(_1300_),
    .X(_0267_));
 sky130_fd_sc_hd__nor2_2 _2689_ (.A(_0881_),
    .B(_0930_),
    .Y(_1301_));
 sky130_fd_sc_hd__mux2_1 _2690_ (.A0(\RAM[67][0] ),
    .A1(_1292_),
    .S(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _2691_ (.A(_1302_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _2692_ (.A0(\RAM[67][1] ),
    .A1(_1295_),
    .S(_1301_),
    .X(_1303_));
 sky130_fd_sc_hd__clkbuf_1 _2693_ (.A(_1303_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(\RAM[67][2] ),
    .A1(_1297_),
    .S(_1301_),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_1 _2695_ (.A(_1304_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _2696_ (.A0(\RAM[67][3] ),
    .A1(_1299_),
    .S(_1301_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_1 _2697_ (.A(_1305_),
    .X(_0271_));
 sky130_fd_sc_hd__nor2_2 _2698_ (.A(_0881_),
    .B(_1039_),
    .Y(_1306_));
 sky130_fd_sc_hd__mux2_1 _2699_ (.A0(\RAM[68][0] ),
    .A1(_1292_),
    .S(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_1 _2700_ (.A(_1307_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _2701_ (.A0(\RAM[68][1] ),
    .A1(_1295_),
    .S(_1306_),
    .X(_1308_));
 sky130_fd_sc_hd__clkbuf_1 _2702_ (.A(_1308_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _2703_ (.A0(\RAM[68][2] ),
    .A1(_1297_),
    .S(_1306_),
    .X(_1309_));
 sky130_fd_sc_hd__clkbuf_1 _2704_ (.A(_1309_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _2705_ (.A0(\RAM[68][3] ),
    .A1(_1299_),
    .S(_1306_),
    .X(_1310_));
 sky130_fd_sc_hd__clkbuf_1 _2706_ (.A(_1310_),
    .X(_0275_));
 sky130_fd_sc_hd__nor2_2 _2707_ (.A(_0978_),
    .B(_1051_),
    .Y(_1311_));
 sky130_fd_sc_hd__mux2_1 _2708_ (.A0(\RAM[6][0] ),
    .A1(_1292_),
    .S(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__clkbuf_1 _2709_ (.A(_1312_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _2710_ (.A0(\RAM[6][1] ),
    .A1(_1295_),
    .S(_1311_),
    .X(_1313_));
 sky130_fd_sc_hd__clkbuf_1 _2711_ (.A(_1313_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _2712_ (.A0(\RAM[6][2] ),
    .A1(_1297_),
    .S(_1311_),
    .X(_1314_));
 sky130_fd_sc_hd__clkbuf_1 _2713_ (.A(_1314_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _2714_ (.A0(\RAM[6][3] ),
    .A1(_1299_),
    .S(_1311_),
    .X(_1315_));
 sky130_fd_sc_hd__clkbuf_1 _2715_ (.A(_1315_),
    .X(_0279_));
 sky130_fd_sc_hd__nor2_2 _2716_ (.A(_0881_),
    .B(_1051_),
    .Y(_1316_));
 sky130_fd_sc_hd__mux2_1 _2717_ (.A0(\RAM[70][0] ),
    .A1(_1292_),
    .S(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__clkbuf_1 _2718_ (.A(_1317_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _2719_ (.A0(\RAM[70][1] ),
    .A1(_1295_),
    .S(_1316_),
    .X(_1318_));
 sky130_fd_sc_hd__clkbuf_1 _2720_ (.A(_1318_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _2721_ (.A0(\RAM[70][2] ),
    .A1(_1297_),
    .S(_1316_),
    .X(_1319_));
 sky130_fd_sc_hd__clkbuf_1 _2722_ (.A(_1319_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _2723_ (.A0(\RAM[70][3] ),
    .A1(_1299_),
    .S(_1316_),
    .X(_1320_));
 sky130_fd_sc_hd__clkbuf_1 _2724_ (.A(_1320_),
    .X(_0283_));
 sky130_fd_sc_hd__nand2_2 _2725_ (.A(_0938_),
    .B(_0922_),
    .Y(_1321_));
 sky130_fd_sc_hd__mux2_1 _2726_ (.A0(_1222_),
    .A1(\RAM[71][0] ),
    .S(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__clkbuf_1 _2727_ (.A(_1322_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _2728_ (.A0(_1226_),
    .A1(\RAM[71][1] ),
    .S(_1321_),
    .X(_1323_));
 sky130_fd_sc_hd__clkbuf_1 _2729_ (.A(_1323_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _2730_ (.A0(_1228_),
    .A1(\RAM[71][2] ),
    .S(_1321_),
    .X(_1324_));
 sky130_fd_sc_hd__clkbuf_1 _2731_ (.A(_1324_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _2732_ (.A0(_1230_),
    .A1(\RAM[71][3] ),
    .S(_1321_),
    .X(_1325_));
 sky130_fd_sc_hd__clkbuf_1 _2733_ (.A(_1325_),
    .X(_0287_));
 sky130_fd_sc_hd__nor2_2 _2734_ (.A(_0881_),
    .B(_1063_),
    .Y(_1326_));
 sky130_fd_sc_hd__mux2_1 _2735_ (.A0(\RAM[72][0] ),
    .A1(_1292_),
    .S(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__clkbuf_1 _2736_ (.A(_1327_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _2737_ (.A0(\RAM[72][1] ),
    .A1(_1295_),
    .S(_1326_),
    .X(_1328_));
 sky130_fd_sc_hd__clkbuf_1 _2738_ (.A(_1328_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _2739_ (.A0(\RAM[72][2] ),
    .A1(_1297_),
    .S(_1326_),
    .X(_1329_));
 sky130_fd_sc_hd__clkbuf_1 _2740_ (.A(_1329_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _2741_ (.A0(\RAM[72][3] ),
    .A1(_1299_),
    .S(_1326_),
    .X(_1330_));
 sky130_fd_sc_hd__clkbuf_1 _2742_ (.A(_1330_),
    .X(_0291_));
 sky130_fd_sc_hd__nor2_2 _2743_ (.A(_0881_),
    .B(_1069_),
    .Y(_1331_));
 sky130_fd_sc_hd__mux2_1 _2744_ (.A0(\RAM[73][0] ),
    .A1(_1292_),
    .S(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_1 _2745_ (.A(_1332_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _2746_ (.A0(\RAM[73][1] ),
    .A1(_1295_),
    .S(_1331_),
    .X(_1333_));
 sky130_fd_sc_hd__clkbuf_1 _2747_ (.A(_1333_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(\RAM[73][2] ),
    .A1(_1297_),
    .S(_1331_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_1 _2749_ (.A(_1334_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _2750_ (.A0(\RAM[73][3] ),
    .A1(_1299_),
    .S(_1331_),
    .X(_1335_));
 sky130_fd_sc_hd__clkbuf_1 _2751_ (.A(_1335_),
    .X(_0295_));
 sky130_fd_sc_hd__nor2_2 _2752_ (.A(_0881_),
    .B(_1076_),
    .Y(_1336_));
 sky130_fd_sc_hd__mux2_1 _2753_ (.A0(\RAM[74][0] ),
    .A1(_1292_),
    .S(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__clkbuf_1 _2754_ (.A(_1337_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _2755_ (.A0(\RAM[74][1] ),
    .A1(_1295_),
    .S(_1336_),
    .X(_1338_));
 sky130_fd_sc_hd__clkbuf_1 _2756_ (.A(_1338_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(\RAM[74][2] ),
    .A1(_1297_),
    .S(_1336_),
    .X(_1339_));
 sky130_fd_sc_hd__clkbuf_1 _2758_ (.A(_1339_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _2759_ (.A0(\RAM[74][3] ),
    .A1(_1299_),
    .S(_1336_),
    .X(_1340_));
 sky130_fd_sc_hd__clkbuf_1 _2760_ (.A(_1340_),
    .X(_0299_));
 sky130_fd_sc_hd__buf_2 _2761_ (.A(_0875_),
    .X(_1341_));
 sky130_fd_sc_hd__nand2_2 _2762_ (.A(_0938_),
    .B(_0905_),
    .Y(_1342_));
 sky130_fd_sc_hd__mux2_1 _2763_ (.A0(_1341_),
    .A1(\RAM[75][0] ),
    .S(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__clkbuf_1 _2764_ (.A(_1343_),
    .X(_0300_));
 sky130_fd_sc_hd__clkbuf_4 _2765_ (.A(_0884_),
    .X(_1344_));
 sky130_fd_sc_hd__mux2_1 _2766_ (.A0(_1344_),
    .A1(\RAM[75][1] ),
    .S(_1342_),
    .X(_1345_));
 sky130_fd_sc_hd__clkbuf_1 _2767_ (.A(_1345_),
    .X(_0301_));
 sky130_fd_sc_hd__buf_2 _2768_ (.A(_0887_),
    .X(_1346_));
 sky130_fd_sc_hd__mux2_1 _2769_ (.A0(_1346_),
    .A1(\RAM[75][2] ),
    .S(_1342_),
    .X(_1347_));
 sky130_fd_sc_hd__clkbuf_1 _2770_ (.A(_1347_),
    .X(_0302_));
 sky130_fd_sc_hd__buf_2 _2771_ (.A(_0890_),
    .X(_1348_));
 sky130_fd_sc_hd__mux2_1 _2772_ (.A0(_1348_),
    .A1(\RAM[75][3] ),
    .S(_1342_),
    .X(_1349_));
 sky130_fd_sc_hd__clkbuf_1 _2773_ (.A(_1349_),
    .X(_0303_));
 sky130_fd_sc_hd__nor2_2 _2774_ (.A(_0880_),
    .B(_0976_),
    .Y(_1350_));
 sky130_fd_sc_hd__mux2_1 _2775_ (.A0(\RAM[76][0] ),
    .A1(_1292_),
    .S(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__clkbuf_1 _2776_ (.A(_1351_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _2777_ (.A0(\RAM[76][1] ),
    .A1(_1295_),
    .S(_1350_),
    .X(_1352_));
 sky130_fd_sc_hd__clkbuf_1 _2778_ (.A(_1352_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _2779_ (.A0(\RAM[76][2] ),
    .A1(_1297_),
    .S(_1350_),
    .X(_1353_));
 sky130_fd_sc_hd__clkbuf_1 _2780_ (.A(_1353_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _2781_ (.A0(\RAM[76][3] ),
    .A1(_1299_),
    .S(_1350_),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_1 _2782_ (.A(_1354_),
    .X(_0307_));
 sky130_fd_sc_hd__nand2_2 _2783_ (.A(_0938_),
    .B(_0946_),
    .Y(_1355_));
 sky130_fd_sc_hd__mux2_1 _2784_ (.A0(_1341_),
    .A1(\RAM[77][0] ),
    .S(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__clkbuf_1 _2785_ (.A(_1356_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _2786_ (.A0(_1344_),
    .A1(\RAM[77][1] ),
    .S(_1355_),
    .X(_1357_));
 sky130_fd_sc_hd__clkbuf_1 _2787_ (.A(_1357_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _2788_ (.A0(_1346_),
    .A1(\RAM[77][2] ),
    .S(_1355_),
    .X(_1358_));
 sky130_fd_sc_hd__clkbuf_1 _2789_ (.A(_1358_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _2790_ (.A0(_1348_),
    .A1(\RAM[77][3] ),
    .S(_1355_),
    .X(_1359_));
 sky130_fd_sc_hd__clkbuf_1 _2791_ (.A(_1359_),
    .X(_0311_));
 sky130_fd_sc_hd__nand2_2 _2792_ (.A(_0938_),
    .B(_0992_),
    .Y(_1360_));
 sky130_fd_sc_hd__mux2_1 _2793_ (.A0(_1341_),
    .A1(\RAM[78][0] ),
    .S(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__clkbuf_1 _2794_ (.A(_1361_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2795_ (.A0(_1344_),
    .A1(\RAM[78][1] ),
    .S(_1360_),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _2796_ (.A(_1362_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2797_ (.A0(_1346_),
    .A1(\RAM[78][2] ),
    .S(_1360_),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_1 _2798_ (.A(_1363_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _2799_ (.A0(_1348_),
    .A1(\RAM[78][3] ),
    .S(_1360_),
    .X(_1364_));
 sky130_fd_sc_hd__clkbuf_1 _2800_ (.A(_1364_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_2 _2801_ (.A(_0922_),
    .B(_0984_),
    .Y(_1365_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(_1341_),
    .A1(\RAM[7][0] ),
    .S(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__clkbuf_1 _2803_ (.A(_1366_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _2804_ (.A0(_1344_),
    .A1(\RAM[7][1] ),
    .S(_1365_),
    .X(_1367_));
 sky130_fd_sc_hd__clkbuf_1 _2805_ (.A(_1367_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _2806_ (.A0(_1346_),
    .A1(\RAM[7][2] ),
    .S(_1365_),
    .X(_1368_));
 sky130_fd_sc_hd__clkbuf_1 _2807_ (.A(_1368_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _2808_ (.A0(_1348_),
    .A1(\RAM[7][3] ),
    .S(_1365_),
    .X(_1369_));
 sky130_fd_sc_hd__clkbuf_1 _2809_ (.A(_1369_),
    .X(_0319_));
 sky130_fd_sc_hd__or2_1 _2810_ (.A(_0601_),
    .B(_0879_),
    .X(_1370_));
 sky130_fd_sc_hd__buf_2 _2811_ (.A(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__nor2_1 _2812_ (.A(_1371_),
    .B(_1007_),
    .Y(_1372_));
 sky130_fd_sc_hd__mux2_1 _2813_ (.A0(\RAM[80][0] ),
    .A1(_1292_),
    .S(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_1 _2814_ (.A(_1373_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _2815_ (.A0(\RAM[80][1] ),
    .A1(_1295_),
    .S(_1372_),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_1 _2816_ (.A(_1374_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _2817_ (.A0(\RAM[80][2] ),
    .A1(_1297_),
    .S(_1372_),
    .X(_1375_));
 sky130_fd_sc_hd__clkbuf_1 _2818_ (.A(_1375_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _2819_ (.A0(\RAM[80][3] ),
    .A1(_1299_),
    .S(_1372_),
    .X(_1376_));
 sky130_fd_sc_hd__clkbuf_1 _2820_ (.A(_1376_),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_4 _2821_ (.A(_0875_),
    .X(_1377_));
 sky130_fd_sc_hd__nor2_2 _2822_ (.A(_1371_),
    .B(_0916_),
    .Y(_1378_));
 sky130_fd_sc_hd__mux2_1 _2823_ (.A0(\RAM[81][0] ),
    .A1(_1377_),
    .S(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _2824_ (.A(_1379_),
    .X(_0324_));
 sky130_fd_sc_hd__buf_4 _2825_ (.A(_0884_),
    .X(_1380_));
 sky130_fd_sc_hd__mux2_1 _2826_ (.A0(\RAM[81][1] ),
    .A1(_1380_),
    .S(_1378_),
    .X(_1381_));
 sky130_fd_sc_hd__clkbuf_1 _2827_ (.A(_1381_),
    .X(_0325_));
 sky130_fd_sc_hd__buf_4 _2828_ (.A(_0887_),
    .X(_1382_));
 sky130_fd_sc_hd__mux2_1 _2829_ (.A0(\RAM[81][2] ),
    .A1(_1382_),
    .S(_1378_),
    .X(_1383_));
 sky130_fd_sc_hd__clkbuf_1 _2830_ (.A(_1383_),
    .X(_0326_));
 sky130_fd_sc_hd__buf_4 _2831_ (.A(_0890_),
    .X(_1384_));
 sky130_fd_sc_hd__mux2_1 _2832_ (.A0(\RAM[81][3] ),
    .A1(_1384_),
    .S(_1378_),
    .X(_1385_));
 sky130_fd_sc_hd__clkbuf_1 _2833_ (.A(_1385_),
    .X(_0327_));
 sky130_fd_sc_hd__nor2_2 _2834_ (.A(_1371_),
    .B(_1021_),
    .Y(_1386_));
 sky130_fd_sc_hd__mux2_1 _2835_ (.A0(\RAM[82][0] ),
    .A1(_1377_),
    .S(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__clkbuf_1 _2836_ (.A(_1387_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _2837_ (.A0(\RAM[82][1] ),
    .A1(_1380_),
    .S(_1386_),
    .X(_1388_));
 sky130_fd_sc_hd__clkbuf_1 _2838_ (.A(_1388_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _2839_ (.A0(\RAM[82][2] ),
    .A1(_1382_),
    .S(_1386_),
    .X(_1389_));
 sky130_fd_sc_hd__clkbuf_1 _2840_ (.A(_1389_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _2841_ (.A0(\RAM[82][3] ),
    .A1(_1384_),
    .S(_1386_),
    .X(_1390_));
 sky130_fd_sc_hd__clkbuf_1 _2842_ (.A(_1390_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_2 _2843_ (.A(_0895_),
    .B(_0952_),
    .Y(_1391_));
 sky130_fd_sc_hd__mux2_1 _2844_ (.A0(_1341_),
    .A1(\RAM[83][0] ),
    .S(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _2845_ (.A(_1392_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _2846_ (.A0(_1344_),
    .A1(\RAM[83][1] ),
    .S(_1391_),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _2847_ (.A(_1393_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _2848_ (.A0(_1346_),
    .A1(\RAM[83][2] ),
    .S(_1391_),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _2849_ (.A(_1394_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _2850_ (.A0(_1348_),
    .A1(\RAM[83][3] ),
    .S(_1391_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_1 _2851_ (.A(_1395_),
    .X(_0335_));
 sky130_fd_sc_hd__nor2_2 _2852_ (.A(_1371_),
    .B(_1039_),
    .Y(_1396_));
 sky130_fd_sc_hd__mux2_1 _2853_ (.A0(\RAM[84][0] ),
    .A1(_1377_),
    .S(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__clkbuf_1 _2854_ (.A(_1397_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _2855_ (.A0(\RAM[84][1] ),
    .A1(_1380_),
    .S(_1396_),
    .X(_1398_));
 sky130_fd_sc_hd__clkbuf_1 _2856_ (.A(_1398_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _2857_ (.A0(\RAM[84][2] ),
    .A1(_1382_),
    .S(_1396_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_1 _2858_ (.A(_1399_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _2859_ (.A0(\RAM[84][3] ),
    .A1(_1384_),
    .S(_1396_),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_1 _2860_ (.A(_1400_),
    .X(_0339_));
 sky130_fd_sc_hd__nand2_2 _2861_ (.A(_1223_),
    .B(_0895_),
    .Y(_1401_));
 sky130_fd_sc_hd__mux2_1 _2862_ (.A0(_1341_),
    .A1(\RAM[85][0] ),
    .S(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__clkbuf_1 _2863_ (.A(_1402_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _2864_ (.A0(_1344_),
    .A1(\RAM[85][1] ),
    .S(_1401_),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_1 _2865_ (.A(_1403_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _2866_ (.A0(_1346_),
    .A1(\RAM[85][2] ),
    .S(_1401_),
    .X(_1404_));
 sky130_fd_sc_hd__clkbuf_1 _2867_ (.A(_1404_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(_1348_),
    .A1(\RAM[85][3] ),
    .S(_1401_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_1 _2869_ (.A(_1405_),
    .X(_0343_));
 sky130_fd_sc_hd__or2_2 _2870_ (.A(_1371_),
    .B(_1051_),
    .X(_1406_));
 sky130_fd_sc_hd__mux2_1 _2871_ (.A0(_1341_),
    .A1(\RAM[86][0] ),
    .S(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__clkbuf_1 _2872_ (.A(_1407_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _2873_ (.A0(_1344_),
    .A1(\RAM[86][1] ),
    .S(_1406_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _2874_ (.A(_1408_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _2875_ (.A0(_1346_),
    .A1(\RAM[86][2] ),
    .S(_1406_),
    .X(_1409_));
 sky130_fd_sc_hd__clkbuf_1 _2876_ (.A(_1409_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _2877_ (.A0(_1348_),
    .A1(\RAM[86][3] ),
    .S(_1406_),
    .X(_1410_));
 sky130_fd_sc_hd__clkbuf_1 _2878_ (.A(_1410_),
    .X(_0347_));
 sky130_fd_sc_hd__nand2_2 _2879_ (.A(_0895_),
    .B(_0922_),
    .Y(_1411_));
 sky130_fd_sc_hd__mux2_1 _2880_ (.A0(_1341_),
    .A1(\RAM[87][0] ),
    .S(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__clkbuf_1 _2881_ (.A(_1412_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _2882_ (.A0(_1344_),
    .A1(\RAM[87][1] ),
    .S(_1411_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_1 _2883_ (.A(_1413_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _2884_ (.A0(_1346_),
    .A1(\RAM[87][2] ),
    .S(_1411_),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _2885_ (.A(_1414_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _2886_ (.A0(_1348_),
    .A1(\RAM[87][3] ),
    .S(_1411_),
    .X(_1415_));
 sky130_fd_sc_hd__clkbuf_1 _2887_ (.A(_1415_),
    .X(_0351_));
 sky130_fd_sc_hd__nor2_2 _2888_ (.A(_1371_),
    .B(_1063_),
    .Y(_1416_));
 sky130_fd_sc_hd__mux2_1 _2889_ (.A0(\RAM[88][0] ),
    .A1(_1377_),
    .S(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__clkbuf_1 _2890_ (.A(_1417_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _2891_ (.A0(\RAM[88][1] ),
    .A1(_1380_),
    .S(_1416_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _2892_ (.A(_1418_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _2893_ (.A0(\RAM[88][2] ),
    .A1(_1382_),
    .S(_1416_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_1 _2894_ (.A(_1419_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _2895_ (.A0(\RAM[88][3] ),
    .A1(_1384_),
    .S(_1416_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _2896_ (.A(_1420_),
    .X(_0355_));
 sky130_fd_sc_hd__nor2_2 _2897_ (.A(_0978_),
    .B(_1063_),
    .Y(_1421_));
 sky130_fd_sc_hd__mux2_1 _2898_ (.A0(\RAM[8][0] ),
    .A1(_1377_),
    .S(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_1 _2899_ (.A(_1422_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _2900_ (.A0(\RAM[8][1] ),
    .A1(_1380_),
    .S(_1421_),
    .X(_1423_));
 sky130_fd_sc_hd__clkbuf_1 _2901_ (.A(_1423_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _2902_ (.A0(\RAM[8][2] ),
    .A1(_1382_),
    .S(_1421_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_1 _2903_ (.A(_1424_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _2904_ (.A0(\RAM[8][3] ),
    .A1(_1384_),
    .S(_1421_),
    .X(_1425_));
 sky130_fd_sc_hd__clkbuf_1 _2905_ (.A(_1425_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_2 _2906_ (.A(_1371_),
    .B(_1076_),
    .X(_1426_));
 sky130_fd_sc_hd__mux2_1 _2907_ (.A0(_1341_),
    .A1(\RAM[90][0] ),
    .S(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__clkbuf_1 _2908_ (.A(_1427_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _2909_ (.A0(_1344_),
    .A1(\RAM[90][1] ),
    .S(_1426_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_1 _2910_ (.A(_1428_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _2911_ (.A0(_1346_),
    .A1(\RAM[90][2] ),
    .S(_1426_),
    .X(_1429_));
 sky130_fd_sc_hd__clkbuf_1 _2912_ (.A(_1429_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _2913_ (.A0(_1348_),
    .A1(\RAM[90][3] ),
    .S(_1426_),
    .X(_1430_));
 sky130_fd_sc_hd__clkbuf_1 _2914_ (.A(_1430_),
    .X(_0363_));
 sky130_fd_sc_hd__nand2_2 _2915_ (.A(_0895_),
    .B(_0905_),
    .Y(_1431_));
 sky130_fd_sc_hd__mux2_1 _2916_ (.A0(_1341_),
    .A1(\RAM[91][0] ),
    .S(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__clkbuf_1 _2917_ (.A(_1432_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _2918_ (.A0(_1344_),
    .A1(\RAM[91][1] ),
    .S(_1431_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _2919_ (.A(_1433_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _2920_ (.A0(_1346_),
    .A1(\RAM[91][2] ),
    .S(_1431_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_1 _2921_ (.A(_1434_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _2922_ (.A0(_1348_),
    .A1(\RAM[91][3] ),
    .S(_1431_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _2923_ (.A(_1435_),
    .X(_0367_));
 sky130_fd_sc_hd__buf_2 _2924_ (.A(_0875_),
    .X(_1436_));
 sky130_fd_sc_hd__or2_2 _2925_ (.A(_1371_),
    .B(_0976_),
    .X(_1437_));
 sky130_fd_sc_hd__mux2_1 _2926_ (.A0(_1436_),
    .A1(\RAM[92][0] ),
    .S(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__clkbuf_1 _2927_ (.A(_1438_),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_4 _2928_ (.A(_0884_),
    .X(_1439_));
 sky130_fd_sc_hd__mux2_1 _2929_ (.A0(_1439_),
    .A1(\RAM[92][1] ),
    .S(_1437_),
    .X(_1440_));
 sky130_fd_sc_hd__clkbuf_1 _2930_ (.A(_1440_),
    .X(_0369_));
 sky130_fd_sc_hd__buf_2 _2931_ (.A(_0887_),
    .X(_1441_));
 sky130_fd_sc_hd__mux2_1 _2932_ (.A0(_1441_),
    .A1(\RAM[92][2] ),
    .S(_1437_),
    .X(_1442_));
 sky130_fd_sc_hd__clkbuf_1 _2933_ (.A(_1442_),
    .X(_0370_));
 sky130_fd_sc_hd__buf_2 _2934_ (.A(_0890_),
    .X(_1443_));
 sky130_fd_sc_hd__mux2_1 _2935_ (.A0(_1443_),
    .A1(\RAM[92][3] ),
    .S(_1437_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _2936_ (.A(_1444_),
    .X(_0371_));
 sky130_fd_sc_hd__nand2_2 _2937_ (.A(_0895_),
    .B(_0946_),
    .Y(_1445_));
 sky130_fd_sc_hd__mux2_1 _2938_ (.A0(_1436_),
    .A1(\RAM[93][0] ),
    .S(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__clkbuf_1 _2939_ (.A(_1446_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _2940_ (.A0(_1439_),
    .A1(\RAM[93][1] ),
    .S(_1445_),
    .X(_1447_));
 sky130_fd_sc_hd__clkbuf_1 _2941_ (.A(_1447_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _2942_ (.A0(_1441_),
    .A1(\RAM[93][2] ),
    .S(_1445_),
    .X(_1448_));
 sky130_fd_sc_hd__clkbuf_1 _2943_ (.A(_1448_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _2944_ (.A0(_1443_),
    .A1(\RAM[93][3] ),
    .S(_1445_),
    .X(_1449_));
 sky130_fd_sc_hd__clkbuf_1 _2945_ (.A(_1449_),
    .X(_0375_));
 sky130_fd_sc_hd__nand2_2 _2946_ (.A(_0895_),
    .B(_0992_),
    .Y(_1450_));
 sky130_fd_sc_hd__mux2_1 _2947_ (.A0(_1436_),
    .A1(\RAM[94][0] ),
    .S(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__clkbuf_1 _2948_ (.A(_1451_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _2949_ (.A0(_1439_),
    .A1(\RAM[94][1] ),
    .S(_1450_),
    .X(_1452_));
 sky130_fd_sc_hd__clkbuf_1 _2950_ (.A(_1452_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _2951_ (.A0(_1441_),
    .A1(\RAM[94][2] ),
    .S(_1450_),
    .X(_1453_));
 sky130_fd_sc_hd__clkbuf_1 _2952_ (.A(_1453_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _2953_ (.A0(_1443_),
    .A1(\RAM[94][3] ),
    .S(_1450_),
    .X(_1454_));
 sky130_fd_sc_hd__clkbuf_1 _2954_ (.A(_1454_),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_2 _2955_ (.A(_0895_),
    .B(_0939_),
    .Y(_1455_));
 sky130_fd_sc_hd__mux2_1 _2956_ (.A0(_1436_),
    .A1(\RAM[95][0] ),
    .S(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__clkbuf_1 _2957_ (.A(_1456_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _2958_ (.A0(_1439_),
    .A1(\RAM[95][1] ),
    .S(_1455_),
    .X(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _2959_ (.A(_1457_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _2960_ (.A0(_1441_),
    .A1(\RAM[95][2] ),
    .S(_1455_),
    .X(_1458_));
 sky130_fd_sc_hd__clkbuf_1 _2961_ (.A(_1458_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _2962_ (.A0(_1443_),
    .A1(\RAM[95][3] ),
    .S(_1455_),
    .X(_1459_));
 sky130_fd_sc_hd__clkbuf_1 _2963_ (.A(_1459_),
    .X(_0383_));
 sky130_fd_sc_hd__or2_1 _2964_ (.A(_0923_),
    .B(_0879_),
    .X(_1460_));
 sky130_fd_sc_hd__clkbuf_4 _2965_ (.A(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__nor2_2 _2966_ (.A(_1461_),
    .B(_1007_),
    .Y(_1462_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(\RAM[96][0] ),
    .A1(_1377_),
    .S(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__clkbuf_1 _2968_ (.A(_1463_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _2969_ (.A0(\RAM[96][1] ),
    .A1(_1380_),
    .S(_1462_),
    .X(_1464_));
 sky130_fd_sc_hd__clkbuf_1 _2970_ (.A(_1464_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _2971_ (.A0(\RAM[96][2] ),
    .A1(_1382_),
    .S(_1462_),
    .X(_1465_));
 sky130_fd_sc_hd__clkbuf_1 _2972_ (.A(_1465_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _2973_ (.A0(\RAM[96][3] ),
    .A1(_1384_),
    .S(_1462_),
    .X(_1466_));
 sky130_fd_sc_hd__clkbuf_1 _2974_ (.A(_1466_),
    .X(_0387_));
 sky130_fd_sc_hd__nor2_2 _2975_ (.A(_0916_),
    .B(_1461_),
    .Y(_1467_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(\RAM[97][0] ),
    .A1(_1377_),
    .S(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _2977_ (.A(_1468_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(\RAM[97][1] ),
    .A1(_1380_),
    .S(_1467_),
    .X(_1469_));
 sky130_fd_sc_hd__clkbuf_1 _2979_ (.A(_1469_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(\RAM[97][2] ),
    .A1(_1382_),
    .S(_1467_),
    .X(_1470_));
 sky130_fd_sc_hd__clkbuf_1 _2981_ (.A(_1470_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(\RAM[97][3] ),
    .A1(_1384_),
    .S(_1467_),
    .X(_1471_));
 sky130_fd_sc_hd__clkbuf_1 _2983_ (.A(_1471_),
    .X(_0391_));
 sky130_fd_sc_hd__nor2_2 _2984_ (.A(_1461_),
    .B(_1021_),
    .Y(_1472_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(\RAM[98][0] ),
    .A1(_1377_),
    .S(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__clkbuf_1 _2986_ (.A(_1473_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _2987_ (.A0(\RAM[98][1] ),
    .A1(_1380_),
    .S(_1472_),
    .X(_1474_));
 sky130_fd_sc_hd__clkbuf_1 _2988_ (.A(_1474_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(\RAM[98][2] ),
    .A1(_1382_),
    .S(_1472_),
    .X(_1475_));
 sky130_fd_sc_hd__clkbuf_1 _2990_ (.A(_1475_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _2991_ (.A0(\RAM[98][3] ),
    .A1(_1384_),
    .S(_1472_),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_1 _2992_ (.A(_1476_),
    .X(_0395_));
 sky130_fd_sc_hd__nor2_2 _2993_ (.A(_0978_),
    .B(_1007_),
    .Y(_1477_));
 sky130_fd_sc_hd__mux2_1 _2994_ (.A0(\RAM[0][0] ),
    .A1(_1377_),
    .S(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_1 _2995_ (.A(_1478_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _2996_ (.A0(\RAM[0][1] ),
    .A1(_1380_),
    .S(_1477_),
    .X(_1479_));
 sky130_fd_sc_hd__clkbuf_1 _2997_ (.A(_1479_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _2998_ (.A0(\RAM[0][2] ),
    .A1(_1382_),
    .S(_1477_),
    .X(_1480_));
 sky130_fd_sc_hd__clkbuf_1 _2999_ (.A(_1480_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _3000_ (.A0(\RAM[0][3] ),
    .A1(_1384_),
    .S(_1477_),
    .X(_1481_));
 sky130_fd_sc_hd__clkbuf_1 _3001_ (.A(_1481_),
    .X(_0399_));
 sky130_fd_sc_hd__nor2_2 _3002_ (.A(_1461_),
    .B(_1039_),
    .Y(_1482_));
 sky130_fd_sc_hd__mux2_1 _3003_ (.A0(\RAM[100][0] ),
    .A1(_1377_),
    .S(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_1 _3004_ (.A(_1483_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _3005_ (.A0(\RAM[100][1] ),
    .A1(_1380_),
    .S(_1482_),
    .X(_1484_));
 sky130_fd_sc_hd__clkbuf_1 _3006_ (.A(_1484_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _3007_ (.A0(\RAM[100][2] ),
    .A1(_1382_),
    .S(_1482_),
    .X(_1485_));
 sky130_fd_sc_hd__clkbuf_1 _3008_ (.A(_1485_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(\RAM[100][3] ),
    .A1(_1384_),
    .S(_1482_),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_1 _3010_ (.A(_1486_),
    .X(_0403_));
 sky130_fd_sc_hd__nand2_2 _3011_ (.A(_1223_),
    .B(_0953_),
    .Y(_1487_));
 sky130_fd_sc_hd__mux2_1 _3012_ (.A0(_1436_),
    .A1(\RAM[101][0] ),
    .S(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__clkbuf_1 _3013_ (.A(_1488_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _3014_ (.A0(_1439_),
    .A1(\RAM[101][1] ),
    .S(_1487_),
    .X(_1489_));
 sky130_fd_sc_hd__clkbuf_1 _3015_ (.A(_1489_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _3016_ (.A0(_1441_),
    .A1(\RAM[101][2] ),
    .S(_1487_),
    .X(_1490_));
 sky130_fd_sc_hd__clkbuf_1 _3017_ (.A(_1490_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(_1443_),
    .A1(\RAM[101][3] ),
    .S(_1487_),
    .X(_1491_));
 sky130_fd_sc_hd__clkbuf_1 _3019_ (.A(_1491_),
    .X(_0407_));
 sky130_fd_sc_hd__or2_2 _3020_ (.A(_1461_),
    .B(_1051_),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_1 _3021_ (.A0(_1436_),
    .A1(\RAM[102][0] ),
    .S(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__clkbuf_1 _3022_ (.A(_1493_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _3023_ (.A0(_1439_),
    .A1(\RAM[102][1] ),
    .S(_1492_),
    .X(_1494_));
 sky130_fd_sc_hd__clkbuf_1 _3024_ (.A(_1494_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _3025_ (.A0(_1441_),
    .A1(\RAM[102][2] ),
    .S(_1492_),
    .X(_1495_));
 sky130_fd_sc_hd__clkbuf_1 _3026_ (.A(_1495_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _3027_ (.A0(_1443_),
    .A1(\RAM[102][3] ),
    .S(_1492_),
    .X(_1496_));
 sky130_fd_sc_hd__clkbuf_1 _3028_ (.A(_1496_),
    .X(_0411_));
 sky130_fd_sc_hd__nand2_2 _3029_ (.A(_0922_),
    .B(_0953_),
    .Y(_1497_));
 sky130_fd_sc_hd__mux2_1 _3030_ (.A0(_1436_),
    .A1(\RAM[103][0] ),
    .S(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__clkbuf_1 _3031_ (.A(_1498_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _3032_ (.A0(_1439_),
    .A1(\RAM[103][1] ),
    .S(_1497_),
    .X(_1499_));
 sky130_fd_sc_hd__clkbuf_1 _3033_ (.A(_1499_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3034_ (.A0(_1441_),
    .A1(\RAM[103][2] ),
    .S(_1497_),
    .X(_1500_));
 sky130_fd_sc_hd__clkbuf_1 _3035_ (.A(_1500_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _3036_ (.A0(_1443_),
    .A1(\RAM[103][3] ),
    .S(_1497_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _3037_ (.A(_1501_),
    .X(_0415_));
 sky130_fd_sc_hd__nor2_2 _3038_ (.A(_1461_),
    .B(_1063_),
    .Y(_1502_));
 sky130_fd_sc_hd__mux2_1 _3039_ (.A0(\RAM[104][0] ),
    .A1(_1018_),
    .S(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__clkbuf_1 _3040_ (.A(_1503_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _3041_ (.A0(\RAM[104][1] ),
    .A1(_1024_),
    .S(_1502_),
    .X(_1504_));
 sky130_fd_sc_hd__clkbuf_1 _3042_ (.A(_1504_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3043_ (.A0(\RAM[104][2] ),
    .A1(_1027_),
    .S(_1502_),
    .X(_1505_));
 sky130_fd_sc_hd__clkbuf_1 _3044_ (.A(_1505_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _3045_ (.A0(\RAM[104][3] ),
    .A1(_1030_),
    .S(_1502_),
    .X(_1506_));
 sky130_fd_sc_hd__clkbuf_1 _3046_ (.A(_1506_),
    .X(_0419_));
 sky130_fd_sc_hd__nand2_2 _3047_ (.A(_0894_),
    .B(_0953_),
    .Y(_1507_));
 sky130_fd_sc_hd__mux2_1 _3048_ (.A0(_1436_),
    .A1(\RAM[105][0] ),
    .S(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__clkbuf_1 _3049_ (.A(_1508_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _3050_ (.A0(_1439_),
    .A1(\RAM[105][1] ),
    .S(_1507_),
    .X(_1509_));
 sky130_fd_sc_hd__clkbuf_1 _3051_ (.A(_1509_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(_1441_),
    .A1(\RAM[105][2] ),
    .S(_1507_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_1 _3053_ (.A(_1510_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _3054_ (.A0(_1443_),
    .A1(\RAM[105][3] ),
    .S(_1507_),
    .X(_1511_));
 sky130_fd_sc_hd__clkbuf_1 _3055_ (.A(_1511_),
    .X(_0423_));
 sky130_fd_sc_hd__or2_2 _3056_ (.A(_1461_),
    .B(_1076_),
    .X(_1512_));
 sky130_fd_sc_hd__mux2_1 _3057_ (.A0(_1436_),
    .A1(\RAM[106][0] ),
    .S(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__clkbuf_1 _3058_ (.A(_1513_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(_1439_),
    .A1(\RAM[106][1] ),
    .S(_1512_),
    .X(_1514_));
 sky130_fd_sc_hd__clkbuf_1 _3060_ (.A(_1514_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(_1441_),
    .A1(\RAM[106][2] ),
    .S(_1512_),
    .X(_1515_));
 sky130_fd_sc_hd__clkbuf_1 _3062_ (.A(_1515_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _3063_ (.A0(_1443_),
    .A1(\RAM[106][3] ),
    .S(_1512_),
    .X(_1516_));
 sky130_fd_sc_hd__clkbuf_1 _3064_ (.A(_1516_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_2 _3065_ (.A(_0905_),
    .B(_0953_),
    .Y(_1517_));
 sky130_fd_sc_hd__mux2_1 _3066_ (.A0(_1436_),
    .A1(\RAM[107][0] ),
    .S(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__clkbuf_1 _3067_ (.A(_1518_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _3068_ (.A0(_1439_),
    .A1(\RAM[107][1] ),
    .S(_1517_),
    .X(_1519_));
 sky130_fd_sc_hd__clkbuf_1 _3069_ (.A(_1519_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _3070_ (.A0(_1441_),
    .A1(\RAM[107][2] ),
    .S(_1517_),
    .X(_1520_));
 sky130_fd_sc_hd__clkbuf_1 _3071_ (.A(_1520_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _3072_ (.A0(_1443_),
    .A1(\RAM[107][3] ),
    .S(_1517_),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_1 _3073_ (.A(_1521_),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_2 _3074_ (.A(_0875_),
    .X(_1522_));
 sky130_fd_sc_hd__or2_2 _3075_ (.A(_1461_),
    .B(_0976_),
    .X(_1523_));
 sky130_fd_sc_hd__mux2_1 _3076_ (.A0(_1522_),
    .A1(\RAM[108][0] ),
    .S(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__clkbuf_1 _3077_ (.A(_1524_),
    .X(_0432_));
 sky130_fd_sc_hd__buf_2 _3078_ (.A(_0884_),
    .X(_1525_));
 sky130_fd_sc_hd__mux2_1 _3079_ (.A0(_1525_),
    .A1(\RAM[108][1] ),
    .S(_1523_),
    .X(_1526_));
 sky130_fd_sc_hd__clkbuf_1 _3080_ (.A(_1526_),
    .X(_0433_));
 sky130_fd_sc_hd__buf_2 _3081_ (.A(_0887_),
    .X(_1527_));
 sky130_fd_sc_hd__mux2_1 _3082_ (.A0(_1527_),
    .A1(\RAM[108][2] ),
    .S(_1523_),
    .X(_1528_));
 sky130_fd_sc_hd__clkbuf_1 _3083_ (.A(_1528_),
    .X(_0434_));
 sky130_fd_sc_hd__buf_2 _3084_ (.A(_0890_),
    .X(_1529_));
 sky130_fd_sc_hd__mux2_1 _3085_ (.A0(_1529_),
    .A1(\RAM[108][3] ),
    .S(_1523_),
    .X(_1530_));
 sky130_fd_sc_hd__clkbuf_1 _3086_ (.A(_1530_),
    .X(_0435_));
 sky130_fd_sc_hd__nor2_2 _3087_ (.A(_0977_),
    .B(_1076_),
    .Y(_1531_));
 sky130_fd_sc_hd__mux2_1 _3088_ (.A0(\RAM[10][0] ),
    .A1(_1018_),
    .S(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_1 _3089_ (.A(_1532_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _3090_ (.A0(\RAM[10][1] ),
    .A1(_1024_),
    .S(_1531_),
    .X(_1533_));
 sky130_fd_sc_hd__clkbuf_1 _3091_ (.A(_1533_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _3092_ (.A0(\RAM[10][2] ),
    .A1(_1027_),
    .S(_1531_),
    .X(_1534_));
 sky130_fd_sc_hd__clkbuf_1 _3093_ (.A(_1534_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _3094_ (.A0(\RAM[10][3] ),
    .A1(_1030_),
    .S(_1531_),
    .X(_1535_));
 sky130_fd_sc_hd__clkbuf_1 _3095_ (.A(_1535_),
    .X(_0439_));
 sky130_fd_sc_hd__nand2_2 _3096_ (.A(_0953_),
    .B(_0992_),
    .Y(_1536_));
 sky130_fd_sc_hd__mux2_1 _3097_ (.A0(_1522_),
    .A1(\RAM[110][0] ),
    .S(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__clkbuf_1 _3098_ (.A(_1537_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _3099_ (.A0(_1525_),
    .A1(\RAM[110][1] ),
    .S(_1536_),
    .X(_1538_));
 sky130_fd_sc_hd__clkbuf_1 _3100_ (.A(_1538_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(_1527_),
    .A1(\RAM[110][2] ),
    .S(_1536_),
    .X(_1539_));
 sky130_fd_sc_hd__clkbuf_1 _3102_ (.A(_1539_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(_1529_),
    .A1(\RAM[110][3] ),
    .S(_1536_),
    .X(_1540_));
 sky130_fd_sc_hd__clkbuf_1 _3104_ (.A(_1540_),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_2 _3105_ (.A(_0939_),
    .B(_0953_),
    .Y(_1541_));
 sky130_fd_sc_hd__mux2_1 _3106_ (.A0(_1522_),
    .A1(\RAM[111][0] ),
    .S(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__clkbuf_1 _3107_ (.A(_1542_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _3108_ (.A0(_1525_),
    .A1(\RAM[111][1] ),
    .S(_1541_),
    .X(_1543_));
 sky130_fd_sc_hd__clkbuf_1 _3109_ (.A(_1543_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _3110_ (.A0(_1527_),
    .A1(\RAM[111][2] ),
    .S(_1541_),
    .X(_1544_));
 sky130_fd_sc_hd__clkbuf_1 _3111_ (.A(_1544_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _3112_ (.A0(_1529_),
    .A1(\RAM[111][3] ),
    .S(_1541_),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_1 _3113_ (.A(_1545_),
    .X(_0447_));
 sky130_fd_sc_hd__or2_1 _3114_ (.A(_0574_),
    .B(_0879_),
    .X(_1546_));
 sky130_fd_sc_hd__clkbuf_4 _3115_ (.A(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__nor2_2 _3116_ (.A(_1547_),
    .B(_1007_),
    .Y(_1548_));
 sky130_fd_sc_hd__mux2_1 _3117_ (.A0(\RAM[112][0] ),
    .A1(_1018_),
    .S(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__clkbuf_1 _3118_ (.A(_1549_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _3119_ (.A0(\RAM[112][1] ),
    .A1(_1024_),
    .S(_1548_),
    .X(_1550_));
 sky130_fd_sc_hd__clkbuf_1 _3120_ (.A(_1550_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _3121_ (.A0(\RAM[112][2] ),
    .A1(_1027_),
    .S(_1548_),
    .X(_1551_));
 sky130_fd_sc_hd__clkbuf_1 _3122_ (.A(_1551_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _3123_ (.A0(\RAM[112][3] ),
    .A1(_1030_),
    .S(_1548_),
    .X(_1552_));
 sky130_fd_sc_hd__clkbuf_1 _3124_ (.A(_1552_),
    .X(_0451_));
 sky130_fd_sc_hd__nor2_2 _3125_ (.A(_0916_),
    .B(_1547_),
    .Y(_1553_));
 sky130_fd_sc_hd__mux2_1 _3126_ (.A0(\RAM[113][0] ),
    .A1(_1018_),
    .S(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__clkbuf_1 _3127_ (.A(_1554_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _3128_ (.A0(\RAM[113][1] ),
    .A1(_1024_),
    .S(_1553_),
    .X(_1555_));
 sky130_fd_sc_hd__clkbuf_1 _3129_ (.A(_1555_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _3130_ (.A0(\RAM[113][2] ),
    .A1(_1027_),
    .S(_1553_),
    .X(_1556_));
 sky130_fd_sc_hd__clkbuf_1 _3131_ (.A(_1556_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _3132_ (.A0(\RAM[113][3] ),
    .A1(_1030_),
    .S(_1553_),
    .X(_1557_));
 sky130_fd_sc_hd__clkbuf_1 _3133_ (.A(_1557_),
    .X(_0455_));
 sky130_fd_sc_hd__nor2_2 _3134_ (.A(_1547_),
    .B(_1021_),
    .Y(_1558_));
 sky130_fd_sc_hd__mux2_1 _3135_ (.A0(\RAM[114][0] ),
    .A1(_1018_),
    .S(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__clkbuf_1 _3136_ (.A(_1559_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _3137_ (.A0(\RAM[114][1] ),
    .A1(_1024_),
    .S(_1558_),
    .X(_1560_));
 sky130_fd_sc_hd__clkbuf_1 _3138_ (.A(_1560_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _3139_ (.A0(\RAM[114][2] ),
    .A1(_1027_),
    .S(_1558_),
    .X(_1561_));
 sky130_fd_sc_hd__clkbuf_1 _3140_ (.A(_1561_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _3141_ (.A0(\RAM[114][3] ),
    .A1(_1030_),
    .S(_1558_),
    .X(_1562_));
 sky130_fd_sc_hd__clkbuf_1 _3142_ (.A(_1562_),
    .X(_0459_));
 sky130_fd_sc_hd__nand2_2 _3143_ (.A(_0952_),
    .B(_0964_),
    .Y(_1563_));
 sky130_fd_sc_hd__mux2_1 _3144_ (.A0(_1522_),
    .A1(\RAM[115][0] ),
    .S(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_1 _3145_ (.A(_1564_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _3146_ (.A0(_1525_),
    .A1(\RAM[115][1] ),
    .S(_1563_),
    .X(_1565_));
 sky130_fd_sc_hd__clkbuf_1 _3147_ (.A(_1565_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _3148_ (.A0(_1527_),
    .A1(\RAM[115][2] ),
    .S(_1563_),
    .X(_1566_));
 sky130_fd_sc_hd__clkbuf_1 _3149_ (.A(_1566_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _3150_ (.A0(_1529_),
    .A1(\RAM[115][3] ),
    .S(_1563_),
    .X(_1567_));
 sky130_fd_sc_hd__clkbuf_1 _3151_ (.A(_1567_),
    .X(_0463_));
 sky130_fd_sc_hd__nor2_2 _3152_ (.A(_1547_),
    .B(_1039_),
    .Y(_1568_));
 sky130_fd_sc_hd__mux2_1 _3153_ (.A0(\RAM[116][0] ),
    .A1(_1018_),
    .S(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__clkbuf_1 _3154_ (.A(_1569_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _3155_ (.A0(\RAM[116][1] ),
    .A1(_1024_),
    .S(_1568_),
    .X(_1570_));
 sky130_fd_sc_hd__clkbuf_1 _3156_ (.A(_1570_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _3157_ (.A0(\RAM[116][2] ),
    .A1(_1027_),
    .S(_1568_),
    .X(_1571_));
 sky130_fd_sc_hd__clkbuf_1 _3158_ (.A(_1571_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _3159_ (.A0(\RAM[116][3] ),
    .A1(_1030_),
    .S(_1568_),
    .X(_1572_));
 sky130_fd_sc_hd__clkbuf_1 _3160_ (.A(_1572_),
    .X(_0467_));
 sky130_fd_sc_hd__nand2_2 _3161_ (.A(_1223_),
    .B(_0964_),
    .Y(_1573_));
 sky130_fd_sc_hd__mux2_1 _3162_ (.A0(_1522_),
    .A1(\RAM[117][0] ),
    .S(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__clkbuf_1 _3163_ (.A(_1574_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _3164_ (.A0(_1525_),
    .A1(\RAM[117][1] ),
    .S(_1573_),
    .X(_1575_));
 sky130_fd_sc_hd__clkbuf_1 _3165_ (.A(_1575_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _3166_ (.A0(_1527_),
    .A1(\RAM[117][2] ),
    .S(_1573_),
    .X(_1576_));
 sky130_fd_sc_hd__clkbuf_1 _3167_ (.A(_1576_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _3168_ (.A0(_1529_),
    .A1(\RAM[117][3] ),
    .S(_1573_),
    .X(_1577_));
 sky130_fd_sc_hd__clkbuf_1 _3169_ (.A(_1577_),
    .X(_0471_));
 sky130_fd_sc_hd__or2_2 _3170_ (.A(_1547_),
    .B(_1051_),
    .X(_1578_));
 sky130_fd_sc_hd__mux2_1 _3171_ (.A0(_1522_),
    .A1(\RAM[118][0] ),
    .S(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__clkbuf_1 _3172_ (.A(_1579_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(_1525_),
    .A1(\RAM[118][1] ),
    .S(_1578_),
    .X(_1580_));
 sky130_fd_sc_hd__clkbuf_1 _3174_ (.A(_1580_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(_1527_),
    .A1(\RAM[118][2] ),
    .S(_1578_),
    .X(_1581_));
 sky130_fd_sc_hd__clkbuf_1 _3176_ (.A(_1581_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _3177_ (.A0(_1529_),
    .A1(\RAM[118][3] ),
    .S(_1578_),
    .X(_1582_));
 sky130_fd_sc_hd__clkbuf_1 _3178_ (.A(_1582_),
    .X(_0475_));
 sky130_fd_sc_hd__nand2_2 _3179_ (.A(_0905_),
    .B(_0984_),
    .Y(_1583_));
 sky130_fd_sc_hd__mux2_1 _3180_ (.A0(_1522_),
    .A1(\RAM[11][0] ),
    .S(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__clkbuf_1 _3181_ (.A(_1584_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _3182_ (.A0(_1525_),
    .A1(\RAM[11][1] ),
    .S(_1583_),
    .X(_1585_));
 sky130_fd_sc_hd__clkbuf_1 _3183_ (.A(_1585_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _3184_ (.A0(_1527_),
    .A1(\RAM[11][2] ),
    .S(_1583_),
    .X(_1586_));
 sky130_fd_sc_hd__clkbuf_1 _3185_ (.A(_1586_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _3186_ (.A0(_1529_),
    .A1(\RAM[11][3] ),
    .S(_1583_),
    .X(_1587_));
 sky130_fd_sc_hd__clkbuf_1 _3187_ (.A(_1587_),
    .X(_0479_));
 sky130_fd_sc_hd__nor2_2 _3188_ (.A(_1547_),
    .B(_1063_),
    .Y(_1588_));
 sky130_fd_sc_hd__mux2_1 _3189_ (.A0(\RAM[120][0] ),
    .A1(_1018_),
    .S(_1588_),
    .X(_1589_));
 sky130_fd_sc_hd__clkbuf_1 _3190_ (.A(_1589_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _3191_ (.A0(\RAM[120][1] ),
    .A1(_1024_),
    .S(_1588_),
    .X(_1590_));
 sky130_fd_sc_hd__clkbuf_1 _3192_ (.A(_1590_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _3193_ (.A0(\RAM[120][2] ),
    .A1(_1027_),
    .S(_1588_),
    .X(_1591_));
 sky130_fd_sc_hd__clkbuf_1 _3194_ (.A(_1591_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _3195_ (.A0(\RAM[120][3] ),
    .A1(_1030_),
    .S(_1588_),
    .X(_1592_));
 sky130_fd_sc_hd__clkbuf_1 _3196_ (.A(_1592_),
    .X(_0483_));
 sky130_fd_sc_hd__nand2_2 _3197_ (.A(_0894_),
    .B(_0964_),
    .Y(_1593_));
 sky130_fd_sc_hd__mux2_1 _3198_ (.A0(_1522_),
    .A1(\RAM[121][0] ),
    .S(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__clkbuf_1 _3199_ (.A(_1594_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(_1525_),
    .A1(\RAM[121][1] ),
    .S(_1593_),
    .X(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _3201_ (.A(_1595_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(_1527_),
    .A1(\RAM[121][2] ),
    .S(_1593_),
    .X(_1596_));
 sky130_fd_sc_hd__clkbuf_1 _3203_ (.A(_1596_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _3204_ (.A0(_1529_),
    .A1(\RAM[121][3] ),
    .S(_1593_),
    .X(_1597_));
 sky130_fd_sc_hd__clkbuf_1 _3205_ (.A(_1597_),
    .X(_0487_));
 sky130_fd_sc_hd__or2_2 _3206_ (.A(_1547_),
    .B(_1076_),
    .X(_1598_));
 sky130_fd_sc_hd__mux2_1 _3207_ (.A0(_1522_),
    .A1(\RAM[122][0] ),
    .S(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__clkbuf_1 _3208_ (.A(_1599_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _3209_ (.A0(_1525_),
    .A1(\RAM[122][1] ),
    .S(_1598_),
    .X(_1600_));
 sky130_fd_sc_hd__clkbuf_1 _3210_ (.A(_1600_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(_1527_),
    .A1(\RAM[122][2] ),
    .S(_1598_),
    .X(_1601_));
 sky130_fd_sc_hd__clkbuf_1 _3212_ (.A(_1601_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _3213_ (.A0(_1529_),
    .A1(\RAM[122][3] ),
    .S(_1598_),
    .X(_1602_));
 sky130_fd_sc_hd__clkbuf_1 _3214_ (.A(_1602_),
    .X(_0491_));
 sky130_fd_sc_hd__nand2_2 _3215_ (.A(_0905_),
    .B(_0964_),
    .Y(_1603_));
 sky130_fd_sc_hd__mux2_1 _3216_ (.A0(_1522_),
    .A1(\RAM[123][0] ),
    .S(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__clkbuf_1 _3217_ (.A(_1604_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(_1525_),
    .A1(\RAM[123][1] ),
    .S(_1603_),
    .X(_1605_));
 sky130_fd_sc_hd__clkbuf_1 _3219_ (.A(_1605_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _3220_ (.A0(_1527_),
    .A1(\RAM[123][2] ),
    .S(_1603_),
    .X(_1606_));
 sky130_fd_sc_hd__clkbuf_1 _3221_ (.A(_1606_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(_1529_),
    .A1(\RAM[123][3] ),
    .S(_1603_),
    .X(_1607_));
 sky130_fd_sc_hd__clkbuf_1 _3223_ (.A(_1607_),
    .X(_0495_));
 sky130_fd_sc_hd__or2_2 _3224_ (.A(_1547_),
    .B(_0976_),
    .X(_1608_));
 sky130_fd_sc_hd__mux2_1 _3225_ (.A0(_0876_),
    .A1(\RAM[124][0] ),
    .S(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__clkbuf_1 _3226_ (.A(_1609_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _3227_ (.A0(_0885_),
    .A1(\RAM[124][1] ),
    .S(_1608_),
    .X(_1610_));
 sky130_fd_sc_hd__clkbuf_1 _3228_ (.A(_1610_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _3229_ (.A0(_0888_),
    .A1(\RAM[124][2] ),
    .S(_1608_),
    .X(_1611_));
 sky130_fd_sc_hd__clkbuf_1 _3230_ (.A(_1611_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _3231_ (.A0(_0891_),
    .A1(\RAM[124][3] ),
    .S(_1608_),
    .X(_1612_));
 sky130_fd_sc_hd__clkbuf_1 _3232_ (.A(_1612_),
    .X(_0499_));
 sky130_fd_sc_hd__nand2_2 _3233_ (.A(_0946_),
    .B(_0964_),
    .Y(_1613_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(_0876_),
    .A1(\RAM[125][0] ),
    .S(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__clkbuf_1 _3235_ (.A(_1614_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _3236_ (.A0(_0885_),
    .A1(\RAM[125][1] ),
    .S(_1613_),
    .X(_1615_));
 sky130_fd_sc_hd__clkbuf_1 _3237_ (.A(_1615_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _3238_ (.A0(_0888_),
    .A1(\RAM[125][2] ),
    .S(_1613_),
    .X(_1616_));
 sky130_fd_sc_hd__clkbuf_1 _3239_ (.A(_1616_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(_0891_),
    .A1(\RAM[125][3] ),
    .S(_1613_),
    .X(_1617_));
 sky130_fd_sc_hd__clkbuf_1 _3241_ (.A(_1617_),
    .X(_0503_));
 sky130_fd_sc_hd__nand2_2 _3242_ (.A(_0964_),
    .B(_0992_),
    .Y(_1618_));
 sky130_fd_sc_hd__mux2_1 _3243_ (.A0(_0876_),
    .A1(\RAM[126][0] ),
    .S(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__clkbuf_1 _3244_ (.A(_1619_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _3245_ (.A0(_0885_),
    .A1(\RAM[126][1] ),
    .S(_1618_),
    .X(_1620_));
 sky130_fd_sc_hd__clkbuf_1 _3246_ (.A(_1620_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _3247_ (.A0(_0888_),
    .A1(\RAM[126][2] ),
    .S(_1618_),
    .X(_1621_));
 sky130_fd_sc_hd__clkbuf_1 _3248_ (.A(_1621_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _3249_ (.A0(_0891_),
    .A1(\RAM[126][3] ),
    .S(_1618_),
    .X(_1622_));
 sky130_fd_sc_hd__clkbuf_1 _3250_ (.A(_1622_),
    .X(_0507_));
 sky130_fd_sc_hd__nor2_2 _3251_ (.A(_1069_),
    .B(_0978_),
    .Y(_1623_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(\RAM[9][0] ),
    .A1(_1018_),
    .S(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__clkbuf_1 _3253_ (.A(_1624_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(\RAM[9][1] ),
    .A1(_1024_),
    .S(_1623_),
    .X(_1625_));
 sky130_fd_sc_hd__clkbuf_1 _3255_ (.A(_1625_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(\RAM[9][2] ),
    .A1(_1027_),
    .S(_1623_),
    .X(_1626_));
 sky130_fd_sc_hd__clkbuf_1 _3257_ (.A(_1626_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(\RAM[9][3] ),
    .A1(_1030_),
    .S(_1623_),
    .X(_1627_));
 sky130_fd_sc_hd__clkbuf_1 _3259_ (.A(_1627_),
    .X(_0511_));
 sky130_fd_sc_hd__dfxtp_1 _3260_ (.CLK(clknet_leaf_24_clk),
    .D(_0000_),
    .Q(\RAM[69][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3261_ (.CLK(clknet_leaf_26_clk),
    .D(_0001_),
    .Q(\RAM[69][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3262_ (.CLK(clknet_leaf_26_clk),
    .D(_0002_),
    .Q(\RAM[69][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3263_ (.CLK(clknet_leaf_26_clk),
    .D(_0003_),
    .Q(\RAM[69][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3264_ (.CLK(clknet_leaf_15_clk),
    .D(_0004_),
    .Q(\RAM[89][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3265_ (.CLK(clknet_leaf_13_clk),
    .D(_0005_),
    .Q(\RAM[89][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3266_ (.CLK(clknet_leaf_14_clk),
    .D(_0006_),
    .Q(\RAM[89][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3267_ (.CLK(clknet_leaf_15_clk),
    .D(_0007_),
    .Q(\RAM[89][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3268_ (.CLK(clknet_leaf_37_clk),
    .D(_0008_),
    .Q(\RAM[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3269_ (.CLK(clknet_leaf_29_clk),
    .D(_0009_),
    .Q(\RAM[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3270_ (.CLK(clknet_leaf_29_clk),
    .D(_0010_),
    .Q(\RAM[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3271_ (.CLK(clknet_leaf_37_clk),
    .D(_0011_),
    .Q(\RAM[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3272_ (.CLK(clknet_leaf_31_clk),
    .D(_0012_),
    .Q(\RAM[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3273_ (.CLK(clknet_leaf_31_clk),
    .D(_0013_),
    .Q(\RAM[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3274_ (.CLK(clknet_leaf_26_clk),
    .D(_0014_),
    .Q(\RAM[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3275_ (.CLK(clknet_leaf_31_clk),
    .D(_0015_),
    .Q(\RAM[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3276_ (.CLK(clknet_leaf_37_clk),
    .D(_0016_),
    .Q(\RAM[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3277_ (.CLK(clknet_leaf_36_clk),
    .D(_0017_),
    .Q(\RAM[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3278_ (.CLK(clknet_leaf_40_clk),
    .D(_0018_),
    .Q(\RAM[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3279_ (.CLK(clknet_leaf_39_clk),
    .D(_0019_),
    .Q(\RAM[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3280_ (.CLK(clknet_leaf_11_clk),
    .D(_0020_),
    .Q(\RAM[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3281_ (.CLK(clknet_leaf_13_clk),
    .D(_0021_),
    .Q(\RAM[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3282_ (.CLK(clknet_leaf_12_clk),
    .D(_0022_),
    .Q(\RAM[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3283_ (.CLK(clknet_leaf_12_clk),
    .D(_0023_),
    .Q(\RAM[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3284_ (.CLK(clknet_leaf_18_clk),
    .D(_0024_),
    .Q(\RAM[79][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3285_ (.CLK(clknet_leaf_20_clk),
    .D(_0025_),
    .Q(\RAM[79][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3286_ (.CLK(clknet_leaf_18_clk),
    .D(_0026_),
    .Q(\RAM[79][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3287_ (.CLK(clknet_leaf_18_clk),
    .D(_0027_),
    .Q(\RAM[79][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3288_ (.CLK(clknet_leaf_11_clk),
    .D(_0028_),
    .Q(\RAM[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3289_ (.CLK(clknet_leaf_11_clk),
    .D(_0029_),
    .Q(\RAM[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3290_ (.CLK(clknet_leaf_6_clk),
    .D(_0030_),
    .Q(\RAM[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3291_ (.CLK(clknet_leaf_11_clk),
    .D(_0031_),
    .Q(\RAM[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3292_ (.CLK(clknet_leaf_0_clk),
    .D(_0032_),
    .Q(\RAM[99][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3293_ (.CLK(clknet_leaf_43_clk),
    .D(_0033_),
    .Q(\RAM[99][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3294_ (.CLK(clknet_leaf_43_clk),
    .D(_0034_),
    .Q(\RAM[99][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3295_ (.CLK(clknet_leaf_43_clk),
    .D(_0035_),
    .Q(\RAM[99][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3296_ (.CLK(clknet_leaf_45_clk),
    .D(_0036_),
    .Q(\RAM[109][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3297_ (.CLK(clknet_leaf_45_clk),
    .D(_0037_),
    .Q(\RAM[109][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3298_ (.CLK(clknet_leaf_43_clk),
    .D(_0038_),
    .Q(\RAM[109][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3299_ (.CLK(clknet_leaf_45_clk),
    .D(_0039_),
    .Q(\RAM[109][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3300_ (.CLK(clknet_leaf_2_clk),
    .D(_0040_),
    .Q(\RAM[119][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3301_ (.CLK(clknet_leaf_1_clk),
    .D(_0041_),
    .Q(\RAM[119][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3302_ (.CLK(clknet_leaf_2_clk),
    .D(_0042_),
    .Q(\RAM[119][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3303_ (.CLK(clknet_leaf_1_clk),
    .D(_0043_),
    .Q(\RAM[119][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3304_ (.CLK(clknet_leaf_38_clk),
    .D(_0044_),
    .Q(\RAM[127][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3305_ (.CLK(clknet_leaf_3_clk),
    .D(_0045_),
    .Q(\RAM[127][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3306_ (.CLK(clknet_leaf_39_clk),
    .D(_0046_),
    .Q(\RAM[127][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3307_ (.CLK(clknet_leaf_39_clk),
    .D(_0047_),
    .Q(\RAM[127][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3308_ (.CLK(clknet_leaf_28_clk),
    .D(_0048_),
    .Q(\RAM[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3309_ (.CLK(clknet_leaf_27_clk),
    .D(_0049_),
    .Q(\RAM[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3310_ (.CLK(clknet_leaf_27_clk),
    .D(_0050_),
    .Q(\RAM[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3311_ (.CLK(clknet_leaf_27_clk),
    .D(_0051_),
    .Q(\RAM[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3312_ (.CLK(clknet_leaf_28_clk),
    .D(_0052_),
    .Q(\RAM[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3313_ (.CLK(clknet_leaf_27_clk),
    .D(_0053_),
    .Q(\RAM[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3314_ (.CLK(clknet_leaf_27_clk),
    .D(_0054_),
    .Q(\RAM[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3315_ (.CLK(clknet_leaf_27_clk),
    .D(_0055_),
    .Q(\RAM[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3316_ (.CLK(clknet_leaf_28_clk),
    .D(_0056_),
    .Q(\RAM[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3317_ (.CLK(clknet_leaf_28_clk),
    .D(_0057_),
    .Q(\RAM[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3318_ (.CLK(clknet_leaf_4_clk),
    .D(_0058_),
    .Q(\RAM[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3319_ (.CLK(clknet_leaf_17_clk),
    .D(_0059_),
    .Q(\RAM[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3320_ (.CLK(clknet_leaf_28_clk),
    .D(_0060_),
    .Q(\RAM[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3321_ (.CLK(clknet_leaf_27_clk),
    .D(_0061_),
    .Q(\RAM[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3322_ (.CLK(clknet_leaf_4_clk),
    .D(_0062_),
    .Q(\RAM[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3323_ (.CLK(clknet_leaf_17_clk),
    .D(_0063_),
    .Q(\RAM[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3324_ (.CLK(clknet_leaf_13_clk),
    .D(_0064_),
    .Q(\RAM[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3325_ (.CLK(clknet_leaf_13_clk),
    .D(_0065_),
    .Q(\RAM[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3326_ (.CLK(clknet_leaf_12_clk),
    .D(_0066_),
    .Q(\RAM[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3327_ (.CLK(clknet_leaf_15_clk),
    .D(_0067_),
    .Q(\RAM[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3328_ (.CLK(clknet_leaf_13_clk),
    .D(_0068_),
    .Q(\RAM[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3329_ (.CLK(clknet_leaf_13_clk),
    .D(_0069_),
    .Q(\RAM[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3330_ (.CLK(clknet_leaf_12_clk),
    .D(_0070_),
    .Q(\RAM[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3331_ (.CLK(clknet_leaf_12_clk),
    .D(_0071_),
    .Q(\RAM[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3332_ (.CLK(clknet_leaf_11_clk),
    .D(_0072_),
    .Q(\RAM[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3333_ (.CLK(clknet_leaf_11_clk),
    .D(_0073_),
    .Q(\RAM[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3334_ (.CLK(clknet_leaf_11_clk),
    .D(_0074_),
    .Q(\RAM[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3335_ (.CLK(clknet_leaf_11_clk),
    .D(_0075_),
    .Q(\RAM[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3336_ (.CLK(clknet_leaf_5_clk),
    .D(_0076_),
    .Q(\RAM[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3337_ (.CLK(clknet_leaf_6_clk),
    .D(_0077_),
    .Q(\RAM[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3338_ (.CLK(clknet_leaf_6_clk),
    .D(_0078_),
    .Q(\RAM[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3339_ (.CLK(clknet_leaf_5_clk),
    .D(_0079_),
    .Q(\RAM[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3340_ (.CLK(clknet_leaf_9_clk),
    .D(_0080_),
    .Q(\RAM[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3341_ (.CLK(clknet_leaf_9_clk),
    .D(_0081_),
    .Q(\RAM[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3342_ (.CLK(clknet_leaf_8_clk),
    .D(_0082_),
    .Q(\RAM[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3343_ (.CLK(clknet_leaf_8_clk),
    .D(_0083_),
    .Q(\RAM[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3344_ (.CLK(clknet_leaf_9_clk),
    .D(_0084_),
    .Q(\RAM[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3345_ (.CLK(clknet_leaf_9_clk),
    .D(_0085_),
    .Q(\RAM[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3346_ (.CLK(clknet_leaf_8_clk),
    .D(_0086_),
    .Q(\RAM[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3347_ (.CLK(clknet_leaf_8_clk),
    .D(_0087_),
    .Q(\RAM[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3348_ (.CLK(clknet_leaf_9_clk),
    .D(_0088_),
    .Q(\RAM[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3349_ (.CLK(clknet_leaf_9_clk),
    .D(_0089_),
    .Q(\RAM[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3350_ (.CLK(clknet_leaf_8_clk),
    .D(_0090_),
    .Q(\RAM[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3351_ (.CLK(clknet_leaf_8_clk),
    .D(_0091_),
    .Q(\RAM[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3352_ (.CLK(clknet_leaf_9_clk),
    .D(_0092_),
    .Q(\RAM[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3353_ (.CLK(clknet_leaf_9_clk),
    .D(_0093_),
    .Q(\RAM[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3354_ (.CLK(clknet_leaf_8_clk),
    .D(_0094_),
    .Q(\RAM[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3355_ (.CLK(clknet_leaf_8_clk),
    .D(_0095_),
    .Q(\RAM[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3356_ (.CLK(clknet_leaf_10_clk),
    .D(_0096_),
    .Q(\RAM[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3357_ (.CLK(clknet_leaf_10_clk),
    .D(_0097_),
    .Q(\RAM[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3358_ (.CLK(clknet_leaf_9_clk),
    .D(_0098_),
    .Q(\RAM[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3359_ (.CLK(clknet_leaf_9_clk),
    .D(_0099_),
    .Q(\RAM[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3360_ (.CLK(clknet_leaf_10_clk),
    .D(_0100_),
    .Q(\RAM[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3361_ (.CLK(clknet_leaf_10_clk),
    .D(_0101_),
    .Q(\RAM[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3362_ (.CLK(clknet_leaf_10_clk),
    .D(_0102_),
    .Q(\RAM[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3363_ (.CLK(clknet_leaf_9_clk),
    .D(_0103_),
    .Q(\RAM[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3364_ (.CLK(clknet_leaf_10_clk),
    .D(_0104_),
    .Q(\RAM[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3365_ (.CLK(clknet_leaf_10_clk),
    .D(_0105_),
    .Q(\RAM[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3366_ (.CLK(clknet_leaf_10_clk),
    .D(_0106_),
    .Q(\RAM[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3367_ (.CLK(clknet_leaf_9_clk),
    .D(_0107_),
    .Q(\RAM[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3368_ (.CLK(clknet_leaf_10_clk),
    .D(_0108_),
    .Q(\RAM[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3369_ (.CLK(clknet_leaf_10_clk),
    .D(_0109_),
    .Q(\RAM[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3370_ (.CLK(clknet_leaf_10_clk),
    .D(_0110_),
    .Q(\RAM[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3371_ (.CLK(clknet_leaf_9_clk),
    .D(_0111_),
    .Q(\RAM[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3372_ (.CLK(clknet_leaf_11_clk),
    .D(_0112_),
    .Q(\RAM[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3373_ (.CLK(clknet_leaf_11_clk),
    .D(_0113_),
    .Q(\RAM[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3374_ (.CLK(clknet_leaf_5_clk),
    .D(_0114_),
    .Q(\RAM[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3375_ (.CLK(clknet_leaf_12_clk),
    .D(_0115_),
    .Q(\RAM[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3376_ (.CLK(clknet_leaf_6_clk),
    .D(_0116_),
    .Q(\RAM[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3377_ (.CLK(clknet_leaf_6_clk),
    .D(_0117_),
    .Q(\RAM[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3378_ (.CLK(clknet_leaf_8_clk),
    .D(_0118_),
    .Q(\RAM[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3379_ (.CLK(clknet_leaf_6_clk),
    .D(_0119_),
    .Q(\RAM[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3380_ (.CLK(clknet_leaf_11_clk),
    .D(_0120_),
    .Q(\RAM[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3381_ (.CLK(clknet_leaf_11_clk),
    .D(_0121_),
    .Q(\RAM[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3382_ (.CLK(clknet_leaf_8_clk),
    .D(_0122_),
    .Q(\RAM[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3383_ (.CLK(clknet_leaf_9_clk),
    .D(_0123_),
    .Q(\RAM[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3384_ (.CLK(clknet_leaf_10_clk),
    .D(_0124_),
    .Q(\RAM[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3385_ (.CLK(clknet_leaf_11_clk),
    .D(_0125_),
    .Q(\RAM[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3386_ (.CLK(clknet_leaf_8_clk),
    .D(_0126_),
    .Q(\RAM[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3387_ (.CLK(clknet_leaf_9_clk),
    .D(_0127_),
    .Q(\RAM[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3388_ (.CLK(clknet_leaf_35_clk),
    .D(_0128_),
    .Q(\RAM[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3389_ (.CLK(clknet_leaf_35_clk),
    .D(_0129_),
    .Q(\RAM[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3390_ (.CLK(clknet_leaf_35_clk),
    .D(_0130_),
    .Q(\RAM[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3391_ (.CLK(clknet_leaf_35_clk),
    .D(_0131_),
    .Q(\RAM[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3392_ (.CLK(clknet_leaf_40_clk),
    .D(_0132_),
    .Q(\RAM[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3393_ (.CLK(clknet_leaf_35_clk),
    .D(_0133_),
    .Q(\RAM[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3394_ (.CLK(clknet_leaf_35_clk),
    .D(_0134_),
    .Q(\RAM[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3395_ (.CLK(clknet_leaf_40_clk),
    .D(_0135_),
    .Q(\RAM[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3396_ (.CLK(clknet_leaf_40_clk),
    .D(_0136_),
    .Q(\RAM[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3397_ (.CLK(clknet_leaf_35_clk),
    .D(_0137_),
    .Q(\RAM[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3398_ (.CLK(clknet_leaf_40_clk),
    .D(_0138_),
    .Q(\RAM[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3399_ (.CLK(clknet_leaf_40_clk),
    .D(_0139_),
    .Q(\RAM[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3400_ (.CLK(clknet_leaf_40_clk),
    .D(_0140_),
    .Q(\RAM[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3401_ (.CLK(clknet_leaf_35_clk),
    .D(_0141_),
    .Q(\RAM[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3402_ (.CLK(clknet_leaf_40_clk),
    .D(_0142_),
    .Q(\RAM[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3403_ (.CLK(clknet_leaf_40_clk),
    .D(_0143_),
    .Q(\RAM[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3404_ (.CLK(clknet_leaf_37_clk),
    .D(_0144_),
    .Q(\RAM[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3405_ (.CLK(clknet_leaf_36_clk),
    .D(_0145_),
    .Q(\RAM[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3406_ (.CLK(clknet_leaf_36_clk),
    .D(_0146_),
    .Q(\RAM[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3407_ (.CLK(clknet_leaf_36_clk),
    .D(_0147_),
    .Q(\RAM[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3408_ (.CLK(clknet_leaf_37_clk),
    .D(_0148_),
    .Q(\RAM[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3409_ (.CLK(clknet_leaf_36_clk),
    .D(_0149_),
    .Q(\RAM[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3410_ (.CLK(clknet_leaf_40_clk),
    .D(_0150_),
    .Q(\RAM[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3411_ (.CLK(clknet_leaf_38_clk),
    .D(_0151_),
    .Q(\RAM[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3412_ (.CLK(clknet_leaf_37_clk),
    .D(_0152_),
    .Q(\RAM[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3413_ (.CLK(clknet_leaf_36_clk),
    .D(_0153_),
    .Q(\RAM[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3414_ (.CLK(clknet_leaf_40_clk),
    .D(_0154_),
    .Q(\RAM[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3415_ (.CLK(clknet_leaf_39_clk),
    .D(_0155_),
    .Q(\RAM[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3416_ (.CLK(clknet_leaf_6_clk),
    .D(_0156_),
    .Q(\RAM[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3417_ (.CLK(clknet_leaf_4_clk),
    .D(_0157_),
    .Q(\RAM[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3418_ (.CLK(clknet_leaf_2_clk),
    .D(_0158_),
    .Q(\RAM[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3419_ (.CLK(clknet_leaf_4_clk),
    .D(_0159_),
    .Q(\RAM[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3420_ (.CLK(clknet_leaf_34_clk),
    .D(_0160_),
    .Q(\RAM[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3421_ (.CLK(clknet_leaf_34_clk),
    .D(_0161_),
    .Q(\RAM[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3422_ (.CLK(clknet_leaf_35_clk),
    .D(_0162_),
    .Q(\RAM[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3423_ (.CLK(clknet_leaf_35_clk),
    .D(_0163_),
    .Q(\RAM[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3424_ (.CLK(clknet_leaf_34_clk),
    .D(_0164_),
    .Q(\RAM[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3425_ (.CLK(clknet_leaf_34_clk),
    .D(_0165_),
    .Q(\RAM[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3426_ (.CLK(clknet_leaf_35_clk),
    .D(_0166_),
    .Q(\RAM[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3427_ (.CLK(clknet_leaf_35_clk),
    .D(_0167_),
    .Q(\RAM[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3428_ (.CLK(clknet_leaf_34_clk),
    .D(_0168_),
    .Q(\RAM[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3429_ (.CLK(clknet_leaf_33_clk),
    .D(_0169_),
    .Q(\RAM[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3430_ (.CLK(clknet_leaf_34_clk),
    .D(_0170_),
    .Q(\RAM[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3431_ (.CLK(clknet_leaf_34_clk),
    .D(_0171_),
    .Q(\RAM[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3432_ (.CLK(clknet_leaf_34_clk),
    .D(_0172_),
    .Q(\RAM[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3433_ (.CLK(clknet_leaf_34_clk),
    .D(_0173_),
    .Q(\RAM[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3434_ (.CLK(clknet_leaf_34_clk),
    .D(_0174_),
    .Q(\RAM[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3435_ (.CLK(clknet_leaf_34_clk),
    .D(_0175_),
    .Q(\RAM[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3436_ (.CLK(clknet_leaf_33_clk),
    .D(_0176_),
    .Q(\RAM[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3437_ (.CLK(clknet_leaf_33_clk),
    .D(_0177_),
    .Q(\RAM[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3438_ (.CLK(clknet_leaf_33_clk),
    .D(_0178_),
    .Q(\RAM[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3439_ (.CLK(clknet_leaf_36_clk),
    .D(_0179_),
    .Q(\RAM[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3440_ (.CLK(clknet_leaf_33_clk),
    .D(_0180_),
    .Q(\RAM[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3441_ (.CLK(clknet_leaf_34_clk),
    .D(_0181_),
    .Q(\RAM[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3442_ (.CLK(clknet_leaf_33_clk),
    .D(_0182_),
    .Q(\RAM[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3443_ (.CLK(clknet_leaf_36_clk),
    .D(_0183_),
    .Q(\RAM[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3444_ (.CLK(clknet_leaf_34_clk),
    .D(_0184_),
    .Q(\RAM[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3445_ (.CLK(clknet_leaf_34_clk),
    .D(_0185_),
    .Q(\RAM[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3446_ (.CLK(clknet_leaf_34_clk),
    .D(_0186_),
    .Q(\RAM[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3447_ (.CLK(clknet_leaf_36_clk),
    .D(_0187_),
    .Q(\RAM[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3448_ (.CLK(clknet_leaf_34_clk),
    .D(_0188_),
    .Q(\RAM[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3449_ (.CLK(clknet_leaf_34_clk),
    .D(_0189_),
    .Q(\RAM[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3450_ (.CLK(clknet_leaf_34_clk),
    .D(_0190_),
    .Q(\RAM[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3451_ (.CLK(clknet_leaf_36_clk),
    .D(_0191_),
    .Q(\RAM[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3452_ (.CLK(clknet_leaf_31_clk),
    .D(_0192_),
    .Q(\RAM[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3453_ (.CLK(clknet_leaf_25_clk),
    .D(_0193_),
    .Q(\RAM[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3454_ (.CLK(clknet_leaf_25_clk),
    .D(_0194_),
    .Q(\RAM[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3455_ (.CLK(clknet_leaf_31_clk),
    .D(_0195_),
    .Q(\RAM[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3456_ (.CLK(clknet_leaf_24_clk),
    .D(_0196_),
    .Q(\RAM[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3457_ (.CLK(clknet_leaf_24_clk),
    .D(_0197_),
    .Q(\RAM[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3458_ (.CLK(clknet_leaf_25_clk),
    .D(_0198_),
    .Q(\RAM[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3459_ (.CLK(clknet_leaf_26_clk),
    .D(_0199_),
    .Q(\RAM[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3460_ (.CLK(clknet_leaf_31_clk),
    .D(_0200_),
    .Q(\RAM[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3461_ (.CLK(clknet_leaf_25_clk),
    .D(_0201_),
    .Q(\RAM[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3462_ (.CLK(clknet_leaf_27_clk),
    .D(_0202_),
    .Q(\RAM[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3463_ (.CLK(clknet_leaf_29_clk),
    .D(_0203_),
    .Q(\RAM[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3464_ (.CLK(clknet_leaf_30_clk),
    .D(_0204_),
    .Q(\RAM[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3465_ (.CLK(clknet_leaf_25_clk),
    .D(_0205_),
    .Q(\RAM[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3466_ (.CLK(clknet_leaf_27_clk),
    .D(_0206_),
    .Q(\RAM[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3467_ (.CLK(clknet_leaf_30_clk),
    .D(_0207_),
    .Q(\RAM[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3468_ (.CLK(clknet_leaf_32_clk),
    .D(_0208_),
    .Q(\RAM[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3469_ (.CLK(clknet_leaf_31_clk),
    .D(_0209_),
    .Q(\RAM[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3470_ (.CLK(clknet_leaf_30_clk),
    .D(_0210_),
    .Q(\RAM[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3471_ (.CLK(clknet_leaf_30_clk),
    .D(_0211_),
    .Q(\RAM[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3472_ (.CLK(clknet_leaf_32_clk),
    .D(_0212_),
    .Q(\RAM[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3473_ (.CLK(clknet_leaf_31_clk),
    .D(_0213_),
    .Q(\RAM[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3474_ (.CLK(clknet_leaf_29_clk),
    .D(_0214_),
    .Q(\RAM[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3475_ (.CLK(clknet_leaf_29_clk),
    .D(_0215_),
    .Q(\RAM[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3476_ (.CLK(clknet_leaf_32_clk),
    .D(_0216_),
    .Q(\RAM[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3477_ (.CLK(clknet_leaf_31_clk),
    .D(_0217_),
    .Q(\RAM[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3478_ (.CLK(clknet_leaf_28_clk),
    .D(_0218_),
    .Q(\RAM[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3479_ (.CLK(clknet_leaf_29_clk),
    .D(_0219_),
    .Q(\RAM[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3480_ (.CLK(clknet_leaf_32_clk),
    .D(_0220_),
    .Q(\RAM[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3481_ (.CLK(clknet_leaf_31_clk),
    .D(_0221_),
    .Q(\RAM[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3482_ (.CLK(clknet_leaf_28_clk),
    .D(_0222_),
    .Q(\RAM[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3483_ (.CLK(clknet_leaf_29_clk),
    .D(_0223_),
    .Q(\RAM[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3484_ (.CLK(clknet_leaf_33_clk),
    .D(_0224_),
    .Q(\RAM[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3485_ (.CLK(clknet_leaf_32_clk),
    .D(_0225_),
    .Q(\RAM[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3486_ (.CLK(clknet_leaf_33_clk),
    .D(_0226_),
    .Q(\RAM[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3487_ (.CLK(clknet_leaf_30_clk),
    .D(_0227_),
    .Q(\RAM[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3488_ (.CLK(clknet_leaf_32_clk),
    .D(_0228_),
    .Q(\RAM[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3489_ (.CLK(clknet_leaf_32_clk),
    .D(_0229_),
    .Q(\RAM[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3490_ (.CLK(clknet_leaf_33_clk),
    .D(_0230_),
    .Q(\RAM[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3491_ (.CLK(clknet_leaf_29_clk),
    .D(_0231_),
    .Q(\RAM[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3492_ (.CLK(clknet_leaf_33_clk),
    .D(_0232_),
    .Q(\RAM[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3493_ (.CLK(clknet_leaf_30_clk),
    .D(_0233_),
    .Q(\RAM[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3494_ (.CLK(clknet_leaf_30_clk),
    .D(_0234_),
    .Q(\RAM[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3495_ (.CLK(clknet_leaf_37_clk),
    .D(_0235_),
    .Q(\RAM[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3496_ (.CLK(clknet_leaf_25_clk),
    .D(_0236_),
    .Q(\RAM[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3497_ (.CLK(clknet_leaf_24_clk),
    .D(_0237_),
    .Q(\RAM[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3498_ (.CLK(clknet_leaf_25_clk),
    .D(_0238_),
    .Q(\RAM[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3499_ (.CLK(clknet_leaf_26_clk),
    .D(_0239_),
    .Q(\RAM[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3500_ (.CLK(clknet_leaf_32_clk),
    .D(_0240_),
    .Q(\RAM[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3501_ (.CLK(clknet_leaf_32_clk),
    .D(_0241_),
    .Q(\RAM[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3502_ (.CLK(clknet_leaf_32_clk),
    .D(_0242_),
    .Q(\RAM[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3503_ (.CLK(clknet_leaf_29_clk),
    .D(_0243_),
    .Q(\RAM[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3504_ (.CLK(clknet_leaf_32_clk),
    .D(_0244_),
    .Q(\RAM[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3505_ (.CLK(clknet_leaf_32_clk),
    .D(_0245_),
    .Q(\RAM[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3506_ (.CLK(clknet_leaf_30_clk),
    .D(_0246_),
    .Q(\RAM[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3507_ (.CLK(clknet_leaf_38_clk),
    .D(_0247_),
    .Q(\RAM[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3508_ (.CLK(clknet_leaf_32_clk),
    .D(_0248_),
    .Q(\RAM[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3509_ (.CLK(clknet_leaf_32_clk),
    .D(_0249_),
    .Q(\RAM[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3510_ (.CLK(clknet_leaf_30_clk),
    .D(_0250_),
    .Q(\RAM[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3511_ (.CLK(clknet_leaf_37_clk),
    .D(_0251_),
    .Q(\RAM[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3512_ (.CLK(clknet_leaf_32_clk),
    .D(_0252_),
    .Q(\RAM[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3513_ (.CLK(clknet_leaf_32_clk),
    .D(_0253_),
    .Q(\RAM[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3514_ (.CLK(clknet_leaf_30_clk),
    .D(_0254_),
    .Q(\RAM[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3515_ (.CLK(clknet_leaf_38_clk),
    .D(_0255_),
    .Q(\RAM[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3516_ (.CLK(clknet_leaf_23_clk),
    .D(_0256_),
    .Q(\RAM[64][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3517_ (.CLK(clknet_leaf_23_clk),
    .D(_0257_),
    .Q(\RAM[64][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3518_ (.CLK(clknet_leaf_23_clk),
    .D(_0258_),
    .Q(\RAM[64][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3519_ (.CLK(clknet_leaf_24_clk),
    .D(_0259_),
    .Q(\RAM[64][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3520_ (.CLK(clknet_leaf_23_clk),
    .D(_0260_),
    .Q(\RAM[65][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3521_ (.CLK(clknet_leaf_23_clk),
    .D(_0261_),
    .Q(\RAM[65][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3522_ (.CLK(clknet_leaf_23_clk),
    .D(_0262_),
    .Q(\RAM[65][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3523_ (.CLK(clknet_leaf_24_clk),
    .D(_0263_),
    .Q(\RAM[65][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3524_ (.CLK(clknet_leaf_23_clk),
    .D(_0264_),
    .Q(\RAM[66][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3525_ (.CLK(clknet_leaf_21_clk),
    .D(_0265_),
    .Q(\RAM[66][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3526_ (.CLK(clknet_leaf_21_clk),
    .D(_0266_),
    .Q(\RAM[66][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3527_ (.CLK(clknet_leaf_23_clk),
    .D(_0267_),
    .Q(\RAM[66][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3528_ (.CLK(clknet_leaf_23_clk),
    .D(_0268_),
    .Q(\RAM[67][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3529_ (.CLK(clknet_leaf_21_clk),
    .D(_0269_),
    .Q(\RAM[67][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3530_ (.CLK(clknet_leaf_23_clk),
    .D(_0270_),
    .Q(\RAM[67][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3531_ (.CLK(clknet_leaf_23_clk),
    .D(_0271_),
    .Q(\RAM[67][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3532_ (.CLK(clknet_leaf_24_clk),
    .D(_0272_),
    .Q(\RAM[68][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3533_ (.CLK(clknet_leaf_24_clk),
    .D(_0273_),
    .Q(\RAM[68][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3534_ (.CLK(clknet_leaf_23_clk),
    .D(_0274_),
    .Q(\RAM[68][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3535_ (.CLK(clknet_leaf_24_clk),
    .D(_0275_),
    .Q(\RAM[68][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3536_ (.CLK(clknet_leaf_27_clk),
    .D(_0276_),
    .Q(\RAM[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3537_ (.CLK(clknet_leaf_17_clk),
    .D(_0277_),
    .Q(\RAM[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3538_ (.CLK(clknet_leaf_27_clk),
    .D(_0278_),
    .Q(\RAM[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3539_ (.CLK(clknet_leaf_17_clk),
    .D(_0279_),
    .Q(\RAM[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3540_ (.CLK(clknet_leaf_24_clk),
    .D(_0280_),
    .Q(\RAM[70][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3541_ (.CLK(clknet_leaf_24_clk),
    .D(_0281_),
    .Q(\RAM[70][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3542_ (.CLK(clknet_leaf_26_clk),
    .D(_0282_),
    .Q(\RAM[70][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3543_ (.CLK(clknet_leaf_26_clk),
    .D(_0283_),
    .Q(\RAM[70][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3544_ (.CLK(clknet_leaf_24_clk),
    .D(_0284_),
    .Q(\RAM[71][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3545_ (.CLK(clknet_leaf_24_clk),
    .D(_0285_),
    .Q(\RAM[71][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3546_ (.CLK(clknet_leaf_26_clk),
    .D(_0286_),
    .Q(\RAM[71][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3547_ (.CLK(clknet_leaf_27_clk),
    .D(_0287_),
    .Q(\RAM[71][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3548_ (.CLK(clknet_leaf_21_clk),
    .D(_0288_),
    .Q(\RAM[72][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3549_ (.CLK(clknet_leaf_22_clk),
    .D(_0289_),
    .Q(\RAM[72][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3550_ (.CLK(clknet_leaf_22_clk),
    .D(_0290_),
    .Q(\RAM[72][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3551_ (.CLK(clknet_leaf_22_clk),
    .D(_0291_),
    .Q(\RAM[72][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3552_ (.CLK(clknet_leaf_21_clk),
    .D(_0292_),
    .Q(\RAM[73][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3553_ (.CLK(clknet_leaf_22_clk),
    .D(_0293_),
    .Q(\RAM[73][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3554_ (.CLK(clknet_leaf_20_clk),
    .D(_0294_),
    .Q(\RAM[73][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3555_ (.CLK(clknet_leaf_22_clk),
    .D(_0295_),
    .Q(\RAM[73][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3556_ (.CLK(clknet_leaf_20_clk),
    .D(_0296_),
    .Q(\RAM[74][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3557_ (.CLK(clknet_leaf_20_clk),
    .D(_0297_),
    .Q(\RAM[74][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3558_ (.CLK(clknet_leaf_20_clk),
    .D(_0298_),
    .Q(\RAM[74][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3559_ (.CLK(clknet_leaf_20_clk),
    .D(_0299_),
    .Q(\RAM[74][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3560_ (.CLK(clknet_leaf_20_clk),
    .D(_0300_),
    .Q(\RAM[75][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3561_ (.CLK(clknet_leaf_20_clk),
    .D(_0301_),
    .Q(\RAM[75][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3562_ (.CLK(clknet_leaf_20_clk),
    .D(_0302_),
    .Q(\RAM[75][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3563_ (.CLK(clknet_leaf_19_clk),
    .D(_0303_),
    .Q(\RAM[75][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3564_ (.CLK(clknet_leaf_21_clk),
    .D(_0304_),
    .Q(\RAM[76][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3565_ (.CLK(clknet_leaf_26_clk),
    .D(_0305_),
    .Q(\RAM[76][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3566_ (.CLK(clknet_leaf_18_clk),
    .D(_0306_),
    .Q(\RAM[76][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3567_ (.CLK(clknet_leaf_18_clk),
    .D(_0307_),
    .Q(\RAM[76][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3568_ (.CLK(clknet_leaf_18_clk),
    .D(_0308_),
    .Q(\RAM[77][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3569_ (.CLK(clknet_leaf_18_clk),
    .D(_0309_),
    .Q(\RAM[77][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3570_ (.CLK(clknet_leaf_18_clk),
    .D(_0310_),
    .Q(\RAM[77][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3571_ (.CLK(clknet_leaf_18_clk),
    .D(_0311_),
    .Q(\RAM[77][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3572_ (.CLK(clknet_leaf_18_clk),
    .D(_0312_),
    .Q(\RAM[78][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3573_ (.CLK(clknet_leaf_20_clk),
    .D(_0313_),
    .Q(\RAM[78][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3574_ (.CLK(clknet_leaf_18_clk),
    .D(_0314_),
    .Q(\RAM[78][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3575_ (.CLK(clknet_leaf_19_clk),
    .D(_0315_),
    .Q(\RAM[78][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3576_ (.CLK(clknet_leaf_27_clk),
    .D(_0316_),
    .Q(\RAM[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3577_ (.CLK(clknet_leaf_16_clk),
    .D(_0317_),
    .Q(\RAM[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3578_ (.CLK(clknet_leaf_27_clk),
    .D(_0318_),
    .Q(\RAM[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3579_ (.CLK(clknet_leaf_17_clk),
    .D(_0319_),
    .Q(\RAM[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3580_ (.CLK(clknet_leaf_18_clk),
    .D(_0320_),
    .Q(\RAM[80][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3581_ (.CLK(clknet_leaf_18_clk),
    .D(_0321_),
    .Q(\RAM[80][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3582_ (.CLK(clknet_leaf_19_clk),
    .D(_0322_),
    .Q(\RAM[80][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3583_ (.CLK(clknet_leaf_19_clk),
    .D(_0323_),
    .Q(\RAM[80][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3584_ (.CLK(clknet_leaf_15_clk),
    .D(_0324_),
    .Q(\RAM[81][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3585_ (.CLK(clknet_leaf_15_clk),
    .D(_0325_),
    .Q(\RAM[81][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3586_ (.CLK(clknet_leaf_14_clk),
    .D(_0326_),
    .Q(\RAM[81][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3587_ (.CLK(clknet_leaf_15_clk),
    .D(_0327_),
    .Q(\RAM[81][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3588_ (.CLK(clknet_leaf_15_clk),
    .D(_0328_),
    .Q(\RAM[82][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3589_ (.CLK(clknet_leaf_15_clk),
    .D(_0329_),
    .Q(\RAM[82][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3590_ (.CLK(clknet_leaf_14_clk),
    .D(_0330_),
    .Q(\RAM[82][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3591_ (.CLK(clknet_leaf_12_clk),
    .D(_0331_),
    .Q(\RAM[82][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3592_ (.CLK(clknet_leaf_16_clk),
    .D(_0332_),
    .Q(\RAM[83][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3593_ (.CLK(clknet_leaf_15_clk),
    .D(_0333_),
    .Q(\RAM[83][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3594_ (.CLK(clknet_leaf_14_clk),
    .D(_0334_),
    .Q(\RAM[83][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3595_ (.CLK(clknet_leaf_12_clk),
    .D(_0335_),
    .Q(\RAM[83][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3596_ (.CLK(clknet_leaf_16_clk),
    .D(_0336_),
    .Q(\RAM[84][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3597_ (.CLK(clknet_leaf_14_clk),
    .D(_0337_),
    .Q(\RAM[84][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3598_ (.CLK(clknet_leaf_19_clk),
    .D(_0338_),
    .Q(\RAM[84][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3599_ (.CLK(clknet_leaf_14_clk),
    .D(_0339_),
    .Q(\RAM[84][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3600_ (.CLK(clknet_leaf_17_clk),
    .D(_0340_),
    .Q(\RAM[85][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3601_ (.CLK(clknet_leaf_20_clk),
    .D(_0341_),
    .Q(\RAM[85][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3602_ (.CLK(clknet_leaf_19_clk),
    .D(_0342_),
    .Q(\RAM[85][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3603_ (.CLK(clknet_leaf_19_clk),
    .D(_0343_),
    .Q(\RAM[85][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3604_ (.CLK(clknet_leaf_17_clk),
    .D(_0344_),
    .Q(\RAM[86][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3605_ (.CLK(clknet_leaf_19_clk),
    .D(_0345_),
    .Q(\RAM[86][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3606_ (.CLK(clknet_leaf_14_clk),
    .D(_0346_),
    .Q(\RAM[86][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3607_ (.CLK(clknet_leaf_19_clk),
    .D(_0347_),
    .Q(\RAM[86][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3608_ (.CLK(clknet_leaf_17_clk),
    .D(_0348_),
    .Q(\RAM[87][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3609_ (.CLK(clknet_leaf_19_clk),
    .D(_0349_),
    .Q(\RAM[87][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3610_ (.CLK(clknet_leaf_19_clk),
    .D(_0350_),
    .Q(\RAM[87][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3611_ (.CLK(clknet_leaf_19_clk),
    .D(_0351_),
    .Q(\RAM[87][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3612_ (.CLK(clknet_leaf_14_clk),
    .D(_0352_),
    .Q(\RAM[88][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3613_ (.CLK(clknet_leaf_13_clk),
    .D(_0353_),
    .Q(\RAM[88][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3614_ (.CLK(clknet_leaf_14_clk),
    .D(_0354_),
    .Q(\RAM[88][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3615_ (.CLK(clknet_leaf_14_clk),
    .D(_0355_),
    .Q(\RAM[88][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3616_ (.CLK(clknet_leaf_6_clk),
    .D(_0356_),
    .Q(\RAM[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3617_ (.CLK(clknet_leaf_7_clk),
    .D(_0357_),
    .Q(\RAM[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3618_ (.CLK(clknet_leaf_6_clk),
    .D(_0358_),
    .Q(\RAM[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3619_ (.CLK(clknet_leaf_7_clk),
    .D(_0359_),
    .Q(\RAM[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3620_ (.CLK(clknet_leaf_15_clk),
    .D(_0360_),
    .Q(\RAM[90][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3621_ (.CLK(clknet_leaf_13_clk),
    .D(_0361_),
    .Q(\RAM[90][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3622_ (.CLK(clknet_leaf_14_clk),
    .D(_0362_),
    .Q(\RAM[90][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3623_ (.CLK(clknet_leaf_13_clk),
    .D(_0363_),
    .Q(\RAM[90][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3624_ (.CLK(clknet_leaf_15_clk),
    .D(_0364_),
    .Q(\RAM[91][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3625_ (.CLK(clknet_leaf_13_clk),
    .D(_0365_),
    .Q(\RAM[91][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3626_ (.CLK(clknet_leaf_14_clk),
    .D(_0366_),
    .Q(\RAM[91][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3627_ (.CLK(clknet_leaf_13_clk),
    .D(_0367_),
    .Q(\RAM[91][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3628_ (.CLK(clknet_leaf_15_clk),
    .D(_0368_),
    .Q(\RAM[92][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3629_ (.CLK(clknet_leaf_4_clk),
    .D(_0369_),
    .Q(\RAM[92][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3630_ (.CLK(clknet_leaf_4_clk),
    .D(_0370_),
    .Q(\RAM[92][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3631_ (.CLK(clknet_leaf_16_clk),
    .D(_0371_),
    .Q(\RAM[92][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3632_ (.CLK(clknet_leaf_16_clk),
    .D(_0372_),
    .Q(\RAM[93][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3633_ (.CLK(clknet_leaf_4_clk),
    .D(_0373_),
    .Q(\RAM[93][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3634_ (.CLK(clknet_leaf_4_clk),
    .D(_0374_),
    .Q(\RAM[93][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3635_ (.CLK(clknet_leaf_4_clk),
    .D(_0375_),
    .Q(\RAM[93][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3636_ (.CLK(clknet_leaf_16_clk),
    .D(_0376_),
    .Q(\RAM[94][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3637_ (.CLK(clknet_leaf_4_clk),
    .D(_0377_),
    .Q(\RAM[94][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3638_ (.CLK(clknet_leaf_4_clk),
    .D(_0378_),
    .Q(\RAM[94][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3639_ (.CLK(clknet_leaf_5_clk),
    .D(_0379_),
    .Q(\RAM[94][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3640_ (.CLK(clknet_leaf_15_clk),
    .D(_0380_),
    .Q(\RAM[95][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3641_ (.CLK(clknet_leaf_4_clk),
    .D(_0381_),
    .Q(\RAM[95][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3642_ (.CLK(clknet_leaf_4_clk),
    .D(_0382_),
    .Q(\RAM[95][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3643_ (.CLK(clknet_leaf_5_clk),
    .D(_0383_),
    .Q(\RAM[95][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3644_ (.CLK(clknet_leaf_39_clk),
    .D(_0384_),
    .Q(\RAM[96][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3645_ (.CLK(clknet_leaf_44_clk),
    .D(_0385_),
    .Q(\RAM[96][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3646_ (.CLK(clknet_leaf_43_clk),
    .D(_0386_),
    .Q(\RAM[96][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3647_ (.CLK(clknet_leaf_42_clk),
    .D(_0387_),
    .Q(\RAM[96][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3648_ (.CLK(clknet_leaf_39_clk),
    .D(_0388_),
    .Q(\RAM[97][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3649_ (.CLK(clknet_leaf_44_clk),
    .D(_0389_),
    .Q(\RAM[97][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3650_ (.CLK(clknet_leaf_45_clk),
    .D(_0390_),
    .Q(\RAM[97][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3651_ (.CLK(clknet_leaf_42_clk),
    .D(_0391_),
    .Q(\RAM[97][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3652_ (.CLK(clknet_leaf_0_clk),
    .D(_0392_),
    .Q(\RAM[98][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3653_ (.CLK(clknet_leaf_44_clk),
    .D(_0393_),
    .Q(\RAM[98][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3654_ (.CLK(clknet_leaf_43_clk),
    .D(_0394_),
    .Q(\RAM[98][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3655_ (.CLK(clknet_leaf_43_clk),
    .D(_0395_),
    .Q(\RAM[98][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3656_ (.CLK(clknet_leaf_5_clk),
    .D(_0396_),
    .Q(\RAM[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3657_ (.CLK(clknet_leaf_5_clk),
    .D(_0397_),
    .Q(\RAM[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3658_ (.CLK(clknet_leaf_6_clk),
    .D(_0398_),
    .Q(\RAM[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3659_ (.CLK(clknet_leaf_5_clk),
    .D(_0399_),
    .Q(\RAM[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3660_ (.CLK(clknet_leaf_39_clk),
    .D(_0400_),
    .Q(\RAM[100][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3661_ (.CLK(clknet_leaf_41_clk),
    .D(_0401_),
    .Q(\RAM[100][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3662_ (.CLK(clknet_leaf_41_clk),
    .D(_0402_),
    .Q(\RAM[100][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3663_ (.CLK(clknet_leaf_40_clk),
    .D(_0403_),
    .Q(\RAM[100][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3664_ (.CLK(clknet_leaf_39_clk),
    .D(_0404_),
    .Q(\RAM[101][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3665_ (.CLK(clknet_leaf_41_clk),
    .D(_0405_),
    .Q(\RAM[101][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3666_ (.CLK(clknet_leaf_41_clk),
    .D(_0406_),
    .Q(\RAM[101][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3667_ (.CLK(clknet_leaf_40_clk),
    .D(_0407_),
    .Q(\RAM[101][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3668_ (.CLK(clknet_leaf_39_clk),
    .D(_0408_),
    .Q(\RAM[102][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3669_ (.CLK(clknet_leaf_41_clk),
    .D(_0409_),
    .Q(\RAM[102][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3670_ (.CLK(clknet_leaf_41_clk),
    .D(_0410_),
    .Q(\RAM[102][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3671_ (.CLK(clknet_leaf_42_clk),
    .D(_0411_),
    .Q(\RAM[102][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3672_ (.CLK(clknet_leaf_39_clk),
    .D(_0412_),
    .Q(\RAM[103][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3673_ (.CLK(clknet_leaf_41_clk),
    .D(_0413_),
    .Q(\RAM[103][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3674_ (.CLK(clknet_leaf_41_clk),
    .D(_0414_),
    .Q(\RAM[103][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3675_ (.CLK(clknet_leaf_42_clk),
    .D(_0415_),
    .Q(\RAM[103][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3676_ (.CLK(clknet_leaf_44_clk),
    .D(_0416_),
    .Q(\RAM[104][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3677_ (.CLK(clknet_leaf_44_clk),
    .D(_0417_),
    .Q(\RAM[104][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3678_ (.CLK(clknet_leaf_44_clk),
    .D(_0418_),
    .Q(\RAM[104][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3679_ (.CLK(clknet_leaf_42_clk),
    .D(_0419_),
    .Q(\RAM[104][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3680_ (.CLK(clknet_leaf_42_clk),
    .D(_0420_),
    .Q(\RAM[105][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3681_ (.CLK(clknet_leaf_44_clk),
    .D(_0421_),
    .Q(\RAM[105][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3682_ (.CLK(clknet_leaf_44_clk),
    .D(_0422_),
    .Q(\RAM[105][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3683_ (.CLK(clknet_leaf_41_clk),
    .D(_0423_),
    .Q(\RAM[105][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3684_ (.CLK(clknet_leaf_42_clk),
    .D(_0424_),
    .Q(\RAM[106][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3685_ (.CLK(clknet_leaf_44_clk),
    .D(_0425_),
    .Q(\RAM[106][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3686_ (.CLK(clknet_leaf_44_clk),
    .D(_0426_),
    .Q(\RAM[106][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3687_ (.CLK(clknet_leaf_42_clk),
    .D(_0427_),
    .Q(\RAM[106][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3688_ (.CLK(clknet_leaf_42_clk),
    .D(_0428_),
    .Q(\RAM[107][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3689_ (.CLK(clknet_leaf_44_clk),
    .D(_0429_),
    .Q(\RAM[107][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3690_ (.CLK(clknet_leaf_44_clk),
    .D(_0430_),
    .Q(\RAM[107][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3691_ (.CLK(clknet_leaf_41_clk),
    .D(_0431_),
    .Q(\RAM[107][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3692_ (.CLK(clknet_leaf_0_clk),
    .D(_0432_),
    .Q(\RAM[108][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3693_ (.CLK(clknet_leaf_45_clk),
    .D(_0433_),
    .Q(\RAM[108][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3694_ (.CLK(clknet_leaf_45_clk),
    .D(_0434_),
    .Q(\RAM[108][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3695_ (.CLK(clknet_leaf_45_clk),
    .D(_0435_),
    .Q(\RAM[108][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3696_ (.CLK(clknet_leaf_6_clk),
    .D(_0436_),
    .Q(\RAM[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3697_ (.CLK(clknet_leaf_7_clk),
    .D(_0437_),
    .Q(\RAM[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3698_ (.CLK(clknet_leaf_7_clk),
    .D(_0438_),
    .Q(\RAM[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3699_ (.CLK(clknet_leaf_7_clk),
    .D(_0439_),
    .Q(\RAM[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3700_ (.CLK(clknet_leaf_45_clk),
    .D(_0440_),
    .Q(\RAM[110][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3701_ (.CLK(clknet_leaf_45_clk),
    .D(_0441_),
    .Q(\RAM[110][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3702_ (.CLK(clknet_leaf_45_clk),
    .D(_0442_),
    .Q(\RAM[110][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3703_ (.CLK(clknet_leaf_45_clk),
    .D(_0443_),
    .Q(\RAM[110][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3704_ (.CLK(clknet_leaf_45_clk),
    .D(_0444_),
    .Q(\RAM[111][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3705_ (.CLK(clknet_leaf_45_clk),
    .D(_0445_),
    .Q(\RAM[111][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3706_ (.CLK(clknet_leaf_45_clk),
    .D(_0446_),
    .Q(\RAM[111][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3707_ (.CLK(clknet_leaf_45_clk),
    .D(_0447_),
    .Q(\RAM[111][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3708_ (.CLK(clknet_leaf_3_clk),
    .D(_0448_),
    .Q(\RAM[112][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3709_ (.CLK(clknet_leaf_3_clk),
    .D(_0449_),
    .Q(\RAM[112][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3710_ (.CLK(clknet_leaf_3_clk),
    .D(_0450_),
    .Q(\RAM[112][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3711_ (.CLK(clknet_leaf_4_clk),
    .D(_0451_),
    .Q(\RAM[112][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3712_ (.CLK(clknet_leaf_3_clk),
    .D(_0452_),
    .Q(\RAM[113][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3713_ (.CLK(clknet_leaf_3_clk),
    .D(_0453_),
    .Q(\RAM[113][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3714_ (.CLK(clknet_leaf_3_clk),
    .D(_0454_),
    .Q(\RAM[113][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3715_ (.CLK(clknet_leaf_4_clk),
    .D(_0455_),
    .Q(\RAM[113][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3716_ (.CLK(clknet_leaf_3_clk),
    .D(_0456_),
    .Q(\RAM[114][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3717_ (.CLK(clknet_leaf_3_clk),
    .D(_0457_),
    .Q(\RAM[114][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3718_ (.CLK(clknet_leaf_3_clk),
    .D(_0458_),
    .Q(\RAM[114][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3719_ (.CLK(clknet_leaf_3_clk),
    .D(_0459_),
    .Q(\RAM[114][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3720_ (.CLK(clknet_leaf_2_clk),
    .D(_0460_),
    .Q(\RAM[115][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3721_ (.CLK(clknet_leaf_3_clk),
    .D(_0461_),
    .Q(\RAM[115][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3722_ (.CLK(clknet_leaf_3_clk),
    .D(_0462_),
    .Q(\RAM[115][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3723_ (.CLK(clknet_leaf_2_clk),
    .D(_0463_),
    .Q(\RAM[115][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3724_ (.CLK(clknet_leaf_2_clk),
    .D(_0464_),
    .Q(\RAM[116][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3725_ (.CLK(clknet_leaf_2_clk),
    .D(_0465_),
    .Q(\RAM[116][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3726_ (.CLK(clknet_leaf_2_clk),
    .D(_0466_),
    .Q(\RAM[116][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3727_ (.CLK(clknet_leaf_1_clk),
    .D(_0467_),
    .Q(\RAM[116][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3728_ (.CLK(clknet_leaf_2_clk),
    .D(_0468_),
    .Q(\RAM[117][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3729_ (.CLK(clknet_leaf_1_clk),
    .D(_0469_),
    .Q(\RAM[117][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3730_ (.CLK(clknet_leaf_3_clk),
    .D(_0470_),
    .Q(\RAM[117][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3731_ (.CLK(clknet_leaf_1_clk),
    .D(_0471_),
    .Q(\RAM[117][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3732_ (.CLK(clknet_leaf_2_clk),
    .D(_0472_),
    .Q(\RAM[118][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3733_ (.CLK(clknet_leaf_1_clk),
    .D(_0473_),
    .Q(\RAM[118][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3734_ (.CLK(clknet_leaf_2_clk),
    .D(_0474_),
    .Q(\RAM[118][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3735_ (.CLK(clknet_leaf_1_clk),
    .D(_0475_),
    .Q(\RAM[118][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3736_ (.CLK(clknet_leaf_6_clk),
    .D(_0476_),
    .Q(\RAM[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3737_ (.CLK(clknet_leaf_7_clk),
    .D(_0477_),
    .Q(\RAM[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3738_ (.CLK(clknet_leaf_6_clk),
    .D(_0478_),
    .Q(\RAM[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3739_ (.CLK(clknet_leaf_7_clk),
    .D(_0479_),
    .Q(\RAM[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3740_ (.CLK(clknet_leaf_3_clk),
    .D(_0480_),
    .Q(\RAM[120][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3741_ (.CLK(clknet_leaf_0_clk),
    .D(_0481_),
    .Q(\RAM[120][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3742_ (.CLK(clknet_leaf_0_clk),
    .D(_0482_),
    .Q(\RAM[120][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3743_ (.CLK(clknet_leaf_0_clk),
    .D(_0483_),
    .Q(\RAM[120][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3744_ (.CLK(clknet_leaf_0_clk),
    .D(_0484_),
    .Q(\RAM[121][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3745_ (.CLK(clknet_leaf_1_clk),
    .D(_0485_),
    .Q(\RAM[121][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3746_ (.CLK(clknet_leaf_0_clk),
    .D(_0486_),
    .Q(\RAM[121][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3747_ (.CLK(clknet_leaf_1_clk),
    .D(_0487_),
    .Q(\RAM[121][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3748_ (.CLK(clknet_leaf_1_clk),
    .D(_0488_),
    .Q(\RAM[122][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3749_ (.CLK(clknet_leaf_1_clk),
    .D(_0489_),
    .Q(\RAM[122][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3750_ (.CLK(clknet_leaf_0_clk),
    .D(_0490_),
    .Q(\RAM[122][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3751_ (.CLK(clknet_leaf_1_clk),
    .D(_0491_),
    .Q(\RAM[122][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3752_ (.CLK(clknet_leaf_1_clk),
    .D(_0492_),
    .Q(\RAM[123][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3753_ (.CLK(clknet_leaf_1_clk),
    .D(_0493_),
    .Q(\RAM[123][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3754_ (.CLK(clknet_leaf_0_clk),
    .D(_0494_),
    .Q(\RAM[123][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3755_ (.CLK(clknet_leaf_1_clk),
    .D(_0495_),
    .Q(\RAM[123][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3756_ (.CLK(clknet_leaf_38_clk),
    .D(_0496_),
    .Q(\RAM[124][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3757_ (.CLK(clknet_leaf_38_clk),
    .D(_0497_),
    .Q(\RAM[124][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3758_ (.CLK(clknet_leaf_38_clk),
    .D(_0498_),
    .Q(\RAM[124][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3759_ (.CLK(clknet_leaf_39_clk),
    .D(_0499_),
    .Q(\RAM[124][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3760_ (.CLK(clknet_leaf_4_clk),
    .D(_0500_),
    .Q(\RAM[125][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3761_ (.CLK(clknet_leaf_38_clk),
    .D(_0501_),
    .Q(\RAM[125][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3762_ (.CLK(clknet_leaf_38_clk),
    .D(_0502_),
    .Q(\RAM[125][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3763_ (.CLK(clknet_leaf_39_clk),
    .D(_0503_),
    .Q(\RAM[125][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3764_ (.CLK(clknet_leaf_4_clk),
    .D(_0504_),
    .Q(\RAM[126][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3765_ (.CLK(clknet_leaf_3_clk),
    .D(_0505_),
    .Q(\RAM[126][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3766_ (.CLK(clknet_leaf_38_clk),
    .D(_0506_),
    .Q(\RAM[126][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3767_ (.CLK(clknet_leaf_3_clk),
    .D(_0507_),
    .Q(\RAM[126][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3768_ (.CLK(clknet_leaf_7_clk),
    .D(_0508_),
    .Q(\RAM[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3769_ (.CLK(clknet_leaf_7_clk),
    .D(_0509_),
    .Q(\RAM[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3770_ (.CLK(clknet_leaf_7_clk),
    .D(_0510_),
    .Q(\RAM[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3771_ (.CLK(clknet_leaf_7_clk),
    .D(_0511_),
    .Q(\RAM[9][3] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(ram_addr[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input2 (.A(ram_addr[1]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(ram_addr[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(ram_addr[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ram_addr[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(ram_addr[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(ram_addr[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(w_val[0]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(w_val[1]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(w_val[2]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(w_val[3]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(wen),
    .X(net12));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(r_val[0]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(r_val[1]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(r_val[2]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(r_val[3]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2145__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2082__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1968__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1954__A1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1842__A1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1805__A1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1670__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1907__C1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__C1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1706__A_N (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1679__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1676__B_N (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1967__A1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__A1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1892__A1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__A1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__A1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1669__A1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1668__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__S1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1971__S1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__S1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__S1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1714__S1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__S1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__S1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1696__A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__S1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__B (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__S1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__S1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1935__S1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__S1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1932__S1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__S1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__S1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1656__S1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1889__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1815__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1663__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1649__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__S0 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1851__S (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1831__S0 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1830__S0 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1828__S0 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1826__S0 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1788__S (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__S0 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1763__S0 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1636__A (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__A (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1822__S0 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__S0 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__S0 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1806__S (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__S0 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1801__S0 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__S0 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1774__S0 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__A (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__A_N (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__S0 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1961__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1955__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1886__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__S0 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__S0 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1658__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__B (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1979__A (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__A (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__A (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__B (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__B (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__B (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__A1 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__A1 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1808__A1 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1793__A1 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1789__A1 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1731__A1 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__A (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1905__S0 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__S0 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1756__S0 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1753__A (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1722__A (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__S (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__A (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__A (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1659__A (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__A (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__S0 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1904__S0 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1901__S0 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__S0 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__S0 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__S0 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1735__S (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__S0 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1678__S0 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__A (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__S0 (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__S (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1850__S (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__S (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__S0 (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1823__S0 (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__S0 (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1733__S (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__S0 (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__S (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1808__B1 (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1789__B1 (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1730__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1647__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1957__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1926__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__C1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__A1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1737__C1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1662__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1648__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__A (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1866__A (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1706__B (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__A (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__A (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__B_N (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1679__A (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1676__A (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1672__A (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__A (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__A1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__A1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1845__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1827__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1790__A1_N (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1757__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1741__A1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1726__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__A1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__A (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__A1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__A (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__A1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__A (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__A1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1796__A1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1668__A1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1657__A (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1978__S (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1976__S (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__S0 (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__S0 (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__S0 (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1765__S0 (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1762__S0 (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1738__A (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__S (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1654__A (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1950__S0 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__S0 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__S0 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__S0 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__S0 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__S0 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1760__S0 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__S0 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__S0 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1655__A (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__S0 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__S (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__S0 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__S0 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1667__S0 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1656__S0 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1989__S0 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__S0 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__S0 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__S0 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__S0 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__S0 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__S0 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__S0 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1712__S0 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1660__A (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2032__A (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__S0 (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1935__S0 (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__S0 (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1932__S0 (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1887__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1812__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1661__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__S1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1831__S1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1830__S1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1828__S1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1826__S1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1763__S1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__A (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1678__S1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1674__A (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1665__A (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__S1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__S1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1852__A (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__S1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1798__S1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1795__S1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1749__S1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__S1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1739__S1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1666__A (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__S1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__S1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__S1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__S1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__A1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1809__A1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__S1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__S1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1732__A1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1667__S1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1670__B (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2104__B (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2070__B (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__B (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1840__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__B2 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__B2 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1692__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__B (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__B (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__B (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__S1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__S1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__S1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1823__S1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__A (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__S1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__S1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__B (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2033__B (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2018__B (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__A1 (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1949__A1 (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__A1 (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1837__A1 (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__B2 (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1764__B2 (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1684__A1 (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2094__B (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2083__B (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__B2 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1949__B2 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__B2 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__A1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1837__B2 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__A1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__A1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1684__B1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__S0 (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__S (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__S (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1786__S (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__S0 (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__A (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1714__S0 (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1710__S0 (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__S0 (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1683__S0 (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__S1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1904__S1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1901__S1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__S1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__S1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__S1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__S1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1710__S1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__S1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1683__S1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__A (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__A (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__A (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1951__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1764__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1691__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__S0 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__S0 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1971__S0 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__S0 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__S0 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__S0 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__S0 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1729__S (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__S0 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__S0 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__A1 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__B1_N (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__A1 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__A1 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__A1 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__B1_N (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1721__A (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__B_N (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1708__A_N (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__A (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2124__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__B1_N (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1951__B1_N (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__B1_N (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__B1_N (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1691__B1_N (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__B2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1981__A1 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1933__B2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1911__B2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__B2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1821__B2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__B2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__B2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__B2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1701__A1 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1981__B2 (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1903__B2 (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1832__B2 (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1750__A (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1716__B2 (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1701__B2 (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1991__A1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__A1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1936__A1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1914__A1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__A1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1824__A1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__A1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__A1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1716__A1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1707__A1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__B2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1903__A1 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1832__A1 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__A1 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1707__B2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1720__C (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1989__S1 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__S1 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__S1 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__S1 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__S1 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__S1 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__S1 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__S1 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__S1 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1712__S1 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__S0 (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__S0 (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__S (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__S0 (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__S0 (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__S (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1780__S0 (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1779__S0 (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__S0 (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1725__S0 (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__S1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__S1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__S1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__S1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__S1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1765__S1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1762__S1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1754__A (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__A (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__A (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__B (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__S1 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1948__S1 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__S1 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__S1 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__S1 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__S1 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1779__S1 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__S1 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1725__S1 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__A (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__A (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__A (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__S0 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__S (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__S0 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__S0 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__S0 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1791__S (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1728__S (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__A (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__B1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1907__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__B1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1829__A (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1814__B1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1793__B1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__S0 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1731__B1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2032__B (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1822__S1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__S1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__S1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1816__S1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__S1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1801__S1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__S1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1774__S1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1925__S (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__S0 (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__S0 (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1816__S0 (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__S0 (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1798__S0 (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1795__S0 (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1749__S0 (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__S0 (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1739__S0 (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__B1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__B1_N (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1833__A1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__A1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__B1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1797__A1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1796__B1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__S1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__C1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1741__B1_N (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1933__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1911__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__B2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1821__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1761__B2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1950__S1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__S1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__S1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__S1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__S1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1780__S1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__S1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1760__S1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__S1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__S1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1991__B2 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__B2 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1936__B2 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1914__B2 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__A1 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__B2 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1824__B2 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__B2 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1761__A1 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__B2 (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__S0 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1987__S0 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__S0 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1948__S0 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1947__S0 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__S0 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1910__S0 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__S0 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__S (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1755__S0 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1987__S1 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__S1 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__A (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__S1 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1947__S1 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__S1 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1910__S1 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__S1 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__S1 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1755__S1 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__D (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__A2 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__B (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__C (.DIODE(_0866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2924__A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2821__A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2166__A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1996__A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__A0 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A0 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A0 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2148__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2050__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2003__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2613__A (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__A (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2249__A (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__A (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__B (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__B (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__B (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2124__B (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__B (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2082__B (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2019__B (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__B (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__A (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2928__A (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2825__A (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__A (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__A (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__A (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__A (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2172__A (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__A (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2006__A (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__A0 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__A0 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A0 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2204__A1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__A1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__A1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__A1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__A1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__A1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__A1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2931__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2010__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__A0 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__A0 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__A0 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__A1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__A1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2186__A1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__A1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2078__A1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2054__A1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__A1 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3084__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2934__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2831__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2686__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2178__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2014__A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__A0 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__A0 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__A0 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2208__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2199__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2154__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2080__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2056__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2158__A0 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2135__A0 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2126__A0 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2116__A0 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2107__A0 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__A0 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__A0 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2062__A0 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2037__A0 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2021__A0 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__A (.DIODE(_0894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__A (.DIODE(_0894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__A (.DIODE(_0894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2020__A (.DIODE(_0894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2160__A0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2137__A0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__A0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2118__A0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__A0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__A0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__A0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__A0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2039__A0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__A0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__A0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2139__A0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2130__A0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2120__A0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__A0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2100__A0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__A0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2066__A0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2041__A0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__A0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2164__A0 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2141__A0 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2132__A0 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__A0 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__A0 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__A0 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__A0 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2068__A0 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2043__A0 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2030__A0 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3179__A (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__A (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2915__B (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__B (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__A (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__A (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__A (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2356__B (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__B (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2145__B (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__B (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2071__B (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2060__B (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__B (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__B (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__A (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2822__B (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__B (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__A (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__A (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2201__A (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2049__B (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3029__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2879__B (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2801__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__B (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__B (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2125__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__A (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2356__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2060__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__B (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__A (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__B (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2073__A (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__A (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__B (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__B (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__B (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2346__B (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2181__A (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2134__A (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__B (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__A (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2937__B (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__B (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__B (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__B (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__A (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2115__A (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2095__B (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__A (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2843__B (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__B (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2106__A (.DIODE(_0952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__B (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__B (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2925__B (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__B (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__B (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__B (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2319__B (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2147__A (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__B (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__A (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2897__A (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__A (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2613__B (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__A (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__B (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__A (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__B (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2147__B (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__A0 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__A0 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__A0 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__A0 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__A0 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2347__A0 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__A0 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__A0 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2270__A0 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2170__A0 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__B (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__B (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__B (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2792__B (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__B (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__B (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__B (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__B (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__A0 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__A0 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__A0 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__A0 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__A0 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__A0 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__A0 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2313__A0 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__A0 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2173__A0 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__A0 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__A0 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__A0 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__A0 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__A0 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__A0 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__A0 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A0 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__A0 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2176__A0 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2543__A0 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__A0 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__A0 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__A0 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__A0 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__A0 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__A0 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__A0 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2276__A0 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2179__A0 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3126__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__A (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__A (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2291__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2261__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2241__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__B (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__B (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2834__B (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2677__B (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__B (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__B (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__B (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__B (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__A1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3137__A1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__A1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__A1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__A1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__A (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__A (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2304__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2293__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2263__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2243__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__A1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__A1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__A1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__A1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__A1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__A1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__A1 (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__A (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__A (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__A1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__A1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2306__A1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2295__A1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__A1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2265__A1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__A1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__A1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__A1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2223__A1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3159__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2367__A (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__A (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__A1 (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__A1 (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__A1 (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__A1 (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__A1 (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__A1 (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__A1 (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__A1 (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__A1 (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2227__A1 (.DIODE(_1031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__B (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__B (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2852__B (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__B (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__B (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__B (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__B (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2240__B (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__B (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__B (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2870__B (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2716__B (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__B (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__B (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__B (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__B (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__B (.DIODE(_1063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__B (.DIODE(_1063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2897__B (.DIODE(_1063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__B (.DIODE(_1063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__B (.DIODE(_1063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__B (.DIODE(_1063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__B (.DIODE(_1063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__B (.DIODE(_1063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__B (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__A (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__A (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3087__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2906__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2301__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2416__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2371__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2400__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2420__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2393__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2422__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2368__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__A1 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__A1 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__A1 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__A1 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__A1 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__A1 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__A1 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__A1 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__A1 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__A1 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__A1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__A1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__A1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__A1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2548__A1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__A1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__A1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__A1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__A1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__A1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__A1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2618__A1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__A1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__A1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__A1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__A1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__A1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__A1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__A1 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__A1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__A1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__A1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__A1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__A1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__A1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__A1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__A1 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2641__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__A0 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__A (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3011__A (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2861__A (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__A (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2643__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2607__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__A0 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__A0 (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2654__A0 (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2645__A0 (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__A0 (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__A0 (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__A0 (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A0 (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__A0 (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__A0 (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__A0 (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__A0 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2656__A0 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__A0 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__A0 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__A0 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__A0 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__A0 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__A0 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__A0 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__A0 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__S (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__S (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__S (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__S (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2813__A1 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__A1 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2753__A1 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__A1 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2735__A1 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__A1 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__A1 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__A1 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__A1 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__A1 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__A1 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__A1 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__A1 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__A1 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__A1 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__A1 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2710__A1 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__A1 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__A1 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2681__A1 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2721__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2694__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2819__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2741__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2723__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2714__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2705__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__S (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__S (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__S (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__S (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__A0 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2907__A0 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__A0 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2871__A0 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2862__A0 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__A0 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__A0 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2793__A0 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__A0 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__A0 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__A0 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2909__A0 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__A0 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2873__A0 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2864__A0 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__A0 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2804__A0 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__A0 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__A0 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__A0 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2920__A0 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2911__A0 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__A0 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2875__A0 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2866__A0 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__A0 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__A0 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2797__A0 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2788__A0 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__A0 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2922__A0 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2913__A0 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2886__A0 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2877__A0 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__A0 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2850__A0 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2808__A0 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__A0 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2790__A0 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__A0 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3003__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2994__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2898__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2889__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2835__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2823__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3005__A1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2996__A1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__A1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__A1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2969__A1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2900__A1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2891__A1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__A1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__A1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__A1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__A1 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2998__A1 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__A1 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__A1 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2971__A1 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2902__A1 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__A1 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2857__A1 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2839__A1 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__A1 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2904__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2895__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2859__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2832__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__A0 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__A0 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3048__A0 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__A0 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3021__A0 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3012__A0 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A0 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__A0 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2938__A0 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2926__A0 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__A0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__A0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__A0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__A0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3023__A0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__A0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__A0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__A0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__A0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2929__A0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__A0 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3061__A0 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__A0 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3034__A0 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__A0 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__A0 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__A0 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__A0 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__A0 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2932__A0 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__A0 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__A0 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__A0 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__A0 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__A0 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__A0 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__A0 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2953__A0 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__A0 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2935__A0 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__A0 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A0 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__A0 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__A0 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__A0 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__A0 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A0 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__A0 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3097__A0 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__A0 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__A0 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__A0 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3200__A0 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__A0 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__A0 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__A0 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__A0 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A0 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__A0 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A0 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__A0 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__A0 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__A0 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__A0 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__A0 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__A0 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__A0 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__A0 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__A0 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3082__A0 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A0 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__A0 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__A0 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A0 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3177__A0 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__A0 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__A0 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__A0 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__A0 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__A0 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__A (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__A (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__A (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__B (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__A (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(ram_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(ram_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(ram_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(ram_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(ram_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(ram_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(ram_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(w_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(w_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(w_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(w_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(wen));
 sky130_fd_sc_hd__diode_2 ANTENNA__1905__S1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__S1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1756__S1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1711__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1664__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1639__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1650__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1672__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__B_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__C1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__C1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1721__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1708__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1628__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__A_N (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1999__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__A1_N (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1843__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1771__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1671__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_output13_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_output14_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_output15_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_output16_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
endmodule

